module chip_top (clk_PAD,
    rst_n_PAD,
    VSS,
    VDD,
    bidir_PAD);
 inout clk_PAD;
 inout rst_n_PAD;
 inout VSS;
 inout VDD;
 inout [53:0] bidir_PAD;

 wire \A_all[0] ;
 wire \A_all[1] ;
 wire \A_all[2] ;
 wire \A_all[3] ;
 wire \A_all[4] ;
 wire \A_all[5] ;
 wire \A_all[6] ;
 wire \A_all[7] ;
 wire \A_all[8] ;
 wire CEN_all;
 wire DAC_clk;
 wire DAC_d1;
 wire DAC_d2;
 wire DAC_le;
 wire \D_all[0] ;
 wire \D_all[1] ;
 wire \D_all[2] ;
 wire \D_all[3] ;
 wire \D_all[4] ;
 wire \D_all[5] ;
 wire \D_all[6] ;
 wire \D_all[7] ;
 wire GWEN_0;
 wire GWEN_1;
 wire GWEN_2;
 wire GWEN_3;
 wire GWEN_4;
 wire GWEN_5;
 wire GWEN_6;
 wire GWEN_7;
 wire \Q0[0] ;
 wire \Q0[1] ;
 wire \Q0[2] ;
 wire \Q0[3] ;
 wire \Q0[4] ;
 wire \Q0[5] ;
 wire \Q0[6] ;
 wire \Q0[7] ;
 wire \Q1[0] ;
 wire \Q1[1] ;
 wire \Q1[2] ;
 wire \Q1[3] ;
 wire \Q1[4] ;
 wire \Q1[5] ;
 wire \Q1[6] ;
 wire \Q1[7] ;
 wire \Q2[0] ;
 wire \Q2[1] ;
 wire \Q2[2] ;
 wire \Q2[3] ;
 wire \Q2[4] ;
 wire \Q2[5] ;
 wire \Q2[6] ;
 wire \Q2[7] ;
 wire \Q3[0] ;
 wire \Q3[1] ;
 wire \Q3[2] ;
 wire \Q3[3] ;
 wire \Q3[4] ;
 wire \Q3[5] ;
 wire \Q3[6] ;
 wire \Q3[7] ;
 wire \Q4[0] ;
 wire \Q4[1] ;
 wire \Q4[2] ;
 wire \Q4[3] ;
 wire \Q4[4] ;
 wire \Q4[5] ;
 wire \Q4[6] ;
 wire \Q4[7] ;
 wire \Q5[0] ;
 wire \Q5[1] ;
 wire \Q5[2] ;
 wire \Q5[3] ;
 wire \Q5[4] ;
 wire \Q5[5] ;
 wire \Q5[6] ;
 wire \Q5[7] ;
 wire \Q6[0] ;
 wire \Q6[1] ;
 wire \Q6[2] ;
 wire \Q6[3] ;
 wire \Q6[4] ;
 wire \Q6[5] ;
 wire \Q6[6] ;
 wire \Q6[7] ;
 wire \Q7[0] ;
 wire \Q7[1] ;
 wire \Q7[2] ;
 wire \Q7[3] ;
 wire \Q7[4] ;
 wire \Q7[5] ;
 wire \Q7[6] ;
 wire \Q7[7] ;
 wire RXD;
 wire TXD;
 wire \WEN_all[0] ;
 wire \WEN_all[1] ;
 wire \WEN_all[2] ;
 wire \WEN_all[3] ;
 wire \WEN_all[4] ;
 wire \WEN_all[5] ;
 wire \WEN_all[6] ;
 wire \WEN_all[7] ;
 wire WEb_ram;
 wire \bidir_CORE2PAD[0] ;
 wire \bidir_CORE2PAD[10] ;
 wire \bidir_CORE2PAD[11] ;
 wire \bidir_CORE2PAD[12] ;
 wire \bidir_CORE2PAD[13] ;
 wire \bidir_CORE2PAD[14] ;
 wire \bidir_CORE2PAD[15] ;
 wire \bidir_CORE2PAD[16] ;
 wire \bidir_CORE2PAD[17] ;
 wire \bidir_CORE2PAD[18] ;
 wire \bidir_CORE2PAD[19] ;
 wire \bidir_CORE2PAD[1] ;
 wire \bidir_CORE2PAD[20] ;
 wire \bidir_CORE2PAD[21] ;
 wire \bidir_CORE2PAD[22] ;
 wire \bidir_CORE2PAD[23] ;
 wire \bidir_CORE2PAD[24] ;
 wire \bidir_CORE2PAD[25] ;
 wire \bidir_CORE2PAD[26] ;
 wire \bidir_CORE2PAD[27] ;
 wire \bidir_CORE2PAD[28] ;
 wire \bidir_CORE2PAD[29] ;
 wire \bidir_CORE2PAD[2] ;
 wire \bidir_CORE2PAD[30] ;
 wire \bidir_CORE2PAD[31] ;
 wire \bidir_CORE2PAD[32] ;
 wire \bidir_CORE2PAD[33] ;
 wire \bidir_CORE2PAD[34] ;
 wire \bidir_CORE2PAD[35] ;
 wire \bidir_CORE2PAD[36] ;
 wire \bidir_CORE2PAD[37] ;
 wire \bidir_CORE2PAD[38] ;
 wire \bidir_CORE2PAD[39] ;
 wire \bidir_CORE2PAD[3] ;
 wire \bidir_CORE2PAD[40] ;
 wire \bidir_CORE2PAD[41] ;
 wire \bidir_CORE2PAD[42] ;
 wire \bidir_CORE2PAD[43] ;
 wire \bidir_CORE2PAD[44] ;
 wire \bidir_CORE2PAD[45] ;
 wire \bidir_CORE2PAD[46] ;
 wire \bidir_CORE2PAD[47] ;
 wire \bidir_CORE2PAD[48] ;
 wire \bidir_CORE2PAD[49] ;
 wire \bidir_CORE2PAD[4] ;
 wire \bidir_CORE2PAD[50] ;
 wire \bidir_CORE2PAD[51] ;
 wire \bidir_CORE2PAD[52] ;
 wire \bidir_CORE2PAD[53] ;
 wire \bidir_CORE2PAD[5] ;
 wire \bidir_CORE2PAD[6] ;
 wire \bidir_CORE2PAD[7] ;
 wire \bidir_CORE2PAD[8] ;
 wire \bidir_CORE2PAD[9] ;
 wire \bidir_CORE2PAD_CS[0] ;
 wire \bidir_CORE2PAD_CS[10] ;
 wire \bidir_CORE2PAD_CS[11] ;
 wire \bidir_CORE2PAD_CS[12] ;
 wire \bidir_CORE2PAD_CS[13] ;
 wire \bidir_CORE2PAD_CS[14] ;
 wire \bidir_CORE2PAD_CS[15] ;
 wire \bidir_CORE2PAD_CS[16] ;
 wire \bidir_CORE2PAD_CS[17] ;
 wire \bidir_CORE2PAD_CS[18] ;
 wire \bidir_CORE2PAD_CS[19] ;
 wire \bidir_CORE2PAD_CS[1] ;
 wire \bidir_CORE2PAD_CS[20] ;
 wire \bidir_CORE2PAD_CS[21] ;
 wire \bidir_CORE2PAD_CS[22] ;
 wire \bidir_CORE2PAD_CS[23] ;
 wire \bidir_CORE2PAD_CS[24] ;
 wire \bidir_CORE2PAD_CS[25] ;
 wire \bidir_CORE2PAD_CS[26] ;
 wire \bidir_CORE2PAD_CS[27] ;
 wire \bidir_CORE2PAD_CS[28] ;
 wire \bidir_CORE2PAD_CS[29] ;
 wire \bidir_CORE2PAD_CS[2] ;
 wire \bidir_CORE2PAD_CS[30] ;
 wire \bidir_CORE2PAD_CS[31] ;
 wire \bidir_CORE2PAD_CS[32] ;
 wire \bidir_CORE2PAD_CS[33] ;
 wire \bidir_CORE2PAD_CS[34] ;
 wire \bidir_CORE2PAD_CS[35] ;
 wire \bidir_CORE2PAD_CS[36] ;
 wire \bidir_CORE2PAD_CS[37] ;
 wire \bidir_CORE2PAD_CS[38] ;
 wire \bidir_CORE2PAD_CS[39] ;
 wire \bidir_CORE2PAD_CS[3] ;
 wire \bidir_CORE2PAD_CS[40] ;
 wire \bidir_CORE2PAD_CS[41] ;
 wire \bidir_CORE2PAD_CS[42] ;
 wire \bidir_CORE2PAD_CS[43] ;
 wire \bidir_CORE2PAD_CS[44] ;
 wire \bidir_CORE2PAD_CS[45] ;
 wire \bidir_CORE2PAD_CS[46] ;
 wire \bidir_CORE2PAD_CS[47] ;
 wire \bidir_CORE2PAD_CS[48] ;
 wire \bidir_CORE2PAD_CS[49] ;
 wire \bidir_CORE2PAD_CS[4] ;
 wire \bidir_CORE2PAD_CS[50] ;
 wire \bidir_CORE2PAD_CS[51] ;
 wire \bidir_CORE2PAD_CS[52] ;
 wire \bidir_CORE2PAD_CS[53] ;
 wire \bidir_CORE2PAD_CS[5] ;
 wire \bidir_CORE2PAD_CS[6] ;
 wire \bidir_CORE2PAD_CS[7] ;
 wire \bidir_CORE2PAD_CS[8] ;
 wire \bidir_CORE2PAD_CS[9] ;
 wire \bidir_CORE2PAD_IE[0] ;
 wire \bidir_CORE2PAD_IE[10] ;
 wire \bidir_CORE2PAD_IE[11] ;
 wire \bidir_CORE2PAD_IE[12] ;
 wire \bidir_CORE2PAD_IE[13] ;
 wire \bidir_CORE2PAD_IE[14] ;
 wire \bidir_CORE2PAD_IE[15] ;
 wire \bidir_CORE2PAD_IE[16] ;
 wire \bidir_CORE2PAD_IE[17] ;
 wire \bidir_CORE2PAD_IE[18] ;
 wire \bidir_CORE2PAD_IE[19] ;
 wire \bidir_CORE2PAD_IE[1] ;
 wire \bidir_CORE2PAD_IE[20] ;
 wire \bidir_CORE2PAD_IE[21] ;
 wire \bidir_CORE2PAD_IE[22] ;
 wire \bidir_CORE2PAD_IE[23] ;
 wire \bidir_CORE2PAD_IE[24] ;
 wire \bidir_CORE2PAD_IE[25] ;
 wire \bidir_CORE2PAD_IE[26] ;
 wire \bidir_CORE2PAD_IE[27] ;
 wire \bidir_CORE2PAD_IE[28] ;
 wire \bidir_CORE2PAD_IE[29] ;
 wire \bidir_CORE2PAD_IE[2] ;
 wire \bidir_CORE2PAD_IE[30] ;
 wire \bidir_CORE2PAD_IE[31] ;
 wire \bidir_CORE2PAD_IE[32] ;
 wire \bidir_CORE2PAD_IE[33] ;
 wire \bidir_CORE2PAD_IE[34] ;
 wire \bidir_CORE2PAD_IE[35] ;
 wire \bidir_CORE2PAD_IE[36] ;
 wire \bidir_CORE2PAD_IE[37] ;
 wire \bidir_CORE2PAD_IE[38] ;
 wire \bidir_CORE2PAD_IE[39] ;
 wire \bidir_CORE2PAD_IE[3] ;
 wire \bidir_CORE2PAD_IE[40] ;
 wire \bidir_CORE2PAD_IE[41] ;
 wire \bidir_CORE2PAD_IE[42] ;
 wire \bidir_CORE2PAD_IE[43] ;
 wire \bidir_CORE2PAD_IE[44] ;
 wire \bidir_CORE2PAD_IE[45] ;
 wire \bidir_CORE2PAD_IE[46] ;
 wire \bidir_CORE2PAD_IE[47] ;
 wire \bidir_CORE2PAD_IE[48] ;
 wire \bidir_CORE2PAD_IE[49] ;
 wire \bidir_CORE2PAD_IE[4] ;
 wire \bidir_CORE2PAD_IE[50] ;
 wire \bidir_CORE2PAD_IE[51] ;
 wire \bidir_CORE2PAD_IE[52] ;
 wire \bidir_CORE2PAD_IE[53] ;
 wire \bidir_CORE2PAD_IE[5] ;
 wire \bidir_CORE2PAD_IE[6] ;
 wire \bidir_CORE2PAD_IE[7] ;
 wire \bidir_CORE2PAD_IE[8] ;
 wire \bidir_CORE2PAD_IE[9] ;
 wire \bidir_CORE2PAD_OE[0] ;
 wire \bidir_CORE2PAD_OE[10] ;
 wire \bidir_CORE2PAD_OE[11] ;
 wire \bidir_CORE2PAD_OE[12] ;
 wire \bidir_CORE2PAD_OE[13] ;
 wire \bidir_CORE2PAD_OE[14] ;
 wire \bidir_CORE2PAD_OE[15] ;
 wire \bidir_CORE2PAD_OE[16] ;
 wire \bidir_CORE2PAD_OE[17] ;
 wire \bidir_CORE2PAD_OE[18] ;
 wire \bidir_CORE2PAD_OE[19] ;
 wire \bidir_CORE2PAD_OE[1] ;
 wire \bidir_CORE2PAD_OE[20] ;
 wire \bidir_CORE2PAD_OE[21] ;
 wire \bidir_CORE2PAD_OE[22] ;
 wire \bidir_CORE2PAD_OE[23] ;
 wire \bidir_CORE2PAD_OE[24] ;
 wire \bidir_CORE2PAD_OE[25] ;
 wire \bidir_CORE2PAD_OE[26] ;
 wire \bidir_CORE2PAD_OE[27] ;
 wire \bidir_CORE2PAD_OE[28] ;
 wire \bidir_CORE2PAD_OE[29] ;
 wire \bidir_CORE2PAD_OE[2] ;
 wire \bidir_CORE2PAD_OE[30] ;
 wire \bidir_CORE2PAD_OE[31] ;
 wire \bidir_CORE2PAD_OE[32] ;
 wire \bidir_CORE2PAD_OE[33] ;
 wire \bidir_CORE2PAD_OE[34] ;
 wire \bidir_CORE2PAD_OE[35] ;
 wire \bidir_CORE2PAD_OE[36] ;
 wire \bidir_CORE2PAD_OE[37] ;
 wire \bidir_CORE2PAD_OE[38] ;
 wire \bidir_CORE2PAD_OE[39] ;
 wire \bidir_CORE2PAD_OE[3] ;
 wire \bidir_CORE2PAD_OE[40] ;
 wire \bidir_CORE2PAD_OE[41] ;
 wire \bidir_CORE2PAD_OE[42] ;
 wire \bidir_CORE2PAD_OE[43] ;
 wire \bidir_CORE2PAD_OE[44] ;
 wire \bidir_CORE2PAD_OE[45] ;
 wire \bidir_CORE2PAD_OE[46] ;
 wire \bidir_CORE2PAD_OE[47] ;
 wire \bidir_CORE2PAD_OE[48] ;
 wire \bidir_CORE2PAD_OE[49] ;
 wire \bidir_CORE2PAD_OE[4] ;
 wire \bidir_CORE2PAD_OE[50] ;
 wire \bidir_CORE2PAD_OE[51] ;
 wire \bidir_CORE2PAD_OE[52] ;
 wire \bidir_CORE2PAD_OE[53] ;
 wire \bidir_CORE2PAD_OE[5] ;
 wire \bidir_CORE2PAD_OE[6] ;
 wire \bidir_CORE2PAD_OE[7] ;
 wire \bidir_CORE2PAD_OE[8] ;
 wire \bidir_CORE2PAD_OE[9] ;
 wire \bidir_CORE2PAD_PD[0] ;
 wire \bidir_CORE2PAD_PD[10] ;
 wire \bidir_CORE2PAD_PD[11] ;
 wire \bidir_CORE2PAD_PD[12] ;
 wire \bidir_CORE2PAD_PD[13] ;
 wire \bidir_CORE2PAD_PD[14] ;
 wire \bidir_CORE2PAD_PD[15] ;
 wire \bidir_CORE2PAD_PD[16] ;
 wire \bidir_CORE2PAD_PD[17] ;
 wire \bidir_CORE2PAD_PD[18] ;
 wire \bidir_CORE2PAD_PD[19] ;
 wire \bidir_CORE2PAD_PD[1] ;
 wire \bidir_CORE2PAD_PD[20] ;
 wire \bidir_CORE2PAD_PD[21] ;
 wire \bidir_CORE2PAD_PD[22] ;
 wire \bidir_CORE2PAD_PD[23] ;
 wire \bidir_CORE2PAD_PD[24] ;
 wire \bidir_CORE2PAD_PD[25] ;
 wire \bidir_CORE2PAD_PD[26] ;
 wire \bidir_CORE2PAD_PD[27] ;
 wire \bidir_CORE2PAD_PD[28] ;
 wire \bidir_CORE2PAD_PD[29] ;
 wire \bidir_CORE2PAD_PD[2] ;
 wire \bidir_CORE2PAD_PD[30] ;
 wire \bidir_CORE2PAD_PD[31] ;
 wire \bidir_CORE2PAD_PD[32] ;
 wire \bidir_CORE2PAD_PD[33] ;
 wire \bidir_CORE2PAD_PD[34] ;
 wire \bidir_CORE2PAD_PD[35] ;
 wire \bidir_CORE2PAD_PD[36] ;
 wire \bidir_CORE2PAD_PD[37] ;
 wire \bidir_CORE2PAD_PD[38] ;
 wire \bidir_CORE2PAD_PD[39] ;
 wire \bidir_CORE2PAD_PD[3] ;
 wire \bidir_CORE2PAD_PD[40] ;
 wire \bidir_CORE2PAD_PD[41] ;
 wire \bidir_CORE2PAD_PD[42] ;
 wire \bidir_CORE2PAD_PD[43] ;
 wire \bidir_CORE2PAD_PD[44] ;
 wire \bidir_CORE2PAD_PD[45] ;
 wire \bidir_CORE2PAD_PD[46] ;
 wire \bidir_CORE2PAD_PD[47] ;
 wire \bidir_CORE2PAD_PD[48] ;
 wire \bidir_CORE2PAD_PD[49] ;
 wire \bidir_CORE2PAD_PD[4] ;
 wire \bidir_CORE2PAD_PD[50] ;
 wire \bidir_CORE2PAD_PD[51] ;
 wire \bidir_CORE2PAD_PD[52] ;
 wire \bidir_CORE2PAD_PD[53] ;
 wire \bidir_CORE2PAD_PD[5] ;
 wire \bidir_CORE2PAD_PD[6] ;
 wire \bidir_CORE2PAD_PD[7] ;
 wire \bidir_CORE2PAD_PD[8] ;
 wire \bidir_CORE2PAD_PD[9] ;
 wire \bidir_CORE2PAD_PU[0] ;
 wire \bidir_CORE2PAD_PU[10] ;
 wire \bidir_CORE2PAD_PU[11] ;
 wire \bidir_CORE2PAD_PU[12] ;
 wire \bidir_CORE2PAD_PU[13] ;
 wire \bidir_CORE2PAD_PU[14] ;
 wire \bidir_CORE2PAD_PU[15] ;
 wire \bidir_CORE2PAD_PU[16] ;
 wire \bidir_CORE2PAD_PU[17] ;
 wire \bidir_CORE2PAD_PU[18] ;
 wire \bidir_CORE2PAD_PU[19] ;
 wire \bidir_CORE2PAD_PU[1] ;
 wire \bidir_CORE2PAD_PU[20] ;
 wire \bidir_CORE2PAD_PU[21] ;
 wire \bidir_CORE2PAD_PU[22] ;
 wire \bidir_CORE2PAD_PU[23] ;
 wire \bidir_CORE2PAD_PU[24] ;
 wire \bidir_CORE2PAD_PU[25] ;
 wire \bidir_CORE2PAD_PU[26] ;
 wire \bidir_CORE2PAD_PU[27] ;
 wire \bidir_CORE2PAD_PU[28] ;
 wire \bidir_CORE2PAD_PU[29] ;
 wire \bidir_CORE2PAD_PU[2] ;
 wire \bidir_CORE2PAD_PU[30] ;
 wire \bidir_CORE2PAD_PU[31] ;
 wire \bidir_CORE2PAD_PU[32] ;
 wire \bidir_CORE2PAD_PU[33] ;
 wire \bidir_CORE2PAD_PU[34] ;
 wire \bidir_CORE2PAD_PU[35] ;
 wire \bidir_CORE2PAD_PU[36] ;
 wire \bidir_CORE2PAD_PU[37] ;
 wire \bidir_CORE2PAD_PU[38] ;
 wire \bidir_CORE2PAD_PU[39] ;
 wire \bidir_CORE2PAD_PU[3] ;
 wire \bidir_CORE2PAD_PU[40] ;
 wire \bidir_CORE2PAD_PU[41] ;
 wire \bidir_CORE2PAD_PU[42] ;
 wire \bidir_CORE2PAD_PU[43] ;
 wire \bidir_CORE2PAD_PU[44] ;
 wire \bidir_CORE2PAD_PU[45] ;
 wire \bidir_CORE2PAD_PU[46] ;
 wire \bidir_CORE2PAD_PU[47] ;
 wire \bidir_CORE2PAD_PU[48] ;
 wire \bidir_CORE2PAD_PU[49] ;
 wire \bidir_CORE2PAD_PU[4] ;
 wire \bidir_CORE2PAD_PU[50] ;
 wire \bidir_CORE2PAD_PU[51] ;
 wire \bidir_CORE2PAD_PU[52] ;
 wire \bidir_CORE2PAD_PU[53] ;
 wire \bidir_CORE2PAD_PU[5] ;
 wire \bidir_CORE2PAD_PU[6] ;
 wire \bidir_CORE2PAD_PU[7] ;
 wire \bidir_CORE2PAD_PU[8] ;
 wire \bidir_CORE2PAD_PU[9] ;
 wire \bidir_CORE2PAD_SL[0] ;
 wire \bidir_CORE2PAD_SL[10] ;
 wire \bidir_CORE2PAD_SL[11] ;
 wire \bidir_CORE2PAD_SL[12] ;
 wire \bidir_CORE2PAD_SL[13] ;
 wire \bidir_CORE2PAD_SL[14] ;
 wire \bidir_CORE2PAD_SL[15] ;
 wire \bidir_CORE2PAD_SL[16] ;
 wire \bidir_CORE2PAD_SL[17] ;
 wire \bidir_CORE2PAD_SL[18] ;
 wire \bidir_CORE2PAD_SL[19] ;
 wire \bidir_CORE2PAD_SL[1] ;
 wire \bidir_CORE2PAD_SL[20] ;
 wire \bidir_CORE2PAD_SL[21] ;
 wire \bidir_CORE2PAD_SL[22] ;
 wire \bidir_CORE2PAD_SL[23] ;
 wire \bidir_CORE2PAD_SL[24] ;
 wire \bidir_CORE2PAD_SL[25] ;
 wire \bidir_CORE2PAD_SL[26] ;
 wire \bidir_CORE2PAD_SL[27] ;
 wire \bidir_CORE2PAD_SL[28] ;
 wire \bidir_CORE2PAD_SL[29] ;
 wire \bidir_CORE2PAD_SL[2] ;
 wire \bidir_CORE2PAD_SL[30] ;
 wire \bidir_CORE2PAD_SL[31] ;
 wire \bidir_CORE2PAD_SL[32] ;
 wire \bidir_CORE2PAD_SL[33] ;
 wire \bidir_CORE2PAD_SL[34] ;
 wire \bidir_CORE2PAD_SL[35] ;
 wire \bidir_CORE2PAD_SL[36] ;
 wire \bidir_CORE2PAD_SL[37] ;
 wire \bidir_CORE2PAD_SL[38] ;
 wire \bidir_CORE2PAD_SL[39] ;
 wire \bidir_CORE2PAD_SL[3] ;
 wire \bidir_CORE2PAD_SL[40] ;
 wire \bidir_CORE2PAD_SL[41] ;
 wire \bidir_CORE2PAD_SL[42] ;
 wire \bidir_CORE2PAD_SL[43] ;
 wire \bidir_CORE2PAD_SL[44] ;
 wire \bidir_CORE2PAD_SL[45] ;
 wire \bidir_CORE2PAD_SL[46] ;
 wire \bidir_CORE2PAD_SL[47] ;
 wire \bidir_CORE2PAD_SL[48] ;
 wire \bidir_CORE2PAD_SL[49] ;
 wire \bidir_CORE2PAD_SL[4] ;
 wire \bidir_CORE2PAD_SL[50] ;
 wire \bidir_CORE2PAD_SL[51] ;
 wire \bidir_CORE2PAD_SL[52] ;
 wire \bidir_CORE2PAD_SL[53] ;
 wire \bidir_CORE2PAD_SL[5] ;
 wire \bidir_CORE2PAD_SL[6] ;
 wire \bidir_CORE2PAD_SL[7] ;
 wire \bidir_CORE2PAD_SL[8] ;
 wire \bidir_CORE2PAD_SL[9] ;
 wire \bidir_PAD2CORE[0] ;
 wire \bidir_PAD2CORE[10] ;
 wire \bidir_PAD2CORE[11] ;
 wire \bidir_PAD2CORE[12] ;
 wire \bidir_PAD2CORE[13] ;
 wire \bidir_PAD2CORE[14] ;
 wire \bidir_PAD2CORE[15] ;
 wire \bidir_PAD2CORE[16] ;
 wire \bidir_PAD2CORE[17] ;
 wire \bidir_PAD2CORE[18] ;
 wire \bidir_PAD2CORE[19] ;
 wire \bidir_PAD2CORE[1] ;
 wire \bidir_PAD2CORE[20] ;
 wire \bidir_PAD2CORE[21] ;
 wire \bidir_PAD2CORE[22] ;
 wire \bidir_PAD2CORE[23] ;
 wire \bidir_PAD2CORE[24] ;
 wire \bidir_PAD2CORE[25] ;
 wire \bidir_PAD2CORE[26] ;
 wire \bidir_PAD2CORE[27] ;
 wire \bidir_PAD2CORE[28] ;
 wire \bidir_PAD2CORE[29] ;
 wire \bidir_PAD2CORE[2] ;
 wire \bidir_PAD2CORE[30] ;
 wire \bidir_PAD2CORE[31] ;
 wire \bidir_PAD2CORE[32] ;
 wire \bidir_PAD2CORE[33] ;
 wire \bidir_PAD2CORE[34] ;
 wire \bidir_PAD2CORE[35] ;
 wire \bidir_PAD2CORE[36] ;
 wire \bidir_PAD2CORE[37] ;
 wire \bidir_PAD2CORE[38] ;
 wire \bidir_PAD2CORE[39] ;
 wire \bidir_PAD2CORE[3] ;
 wire \bidir_PAD2CORE[40] ;
 wire \bidir_PAD2CORE[41] ;
 wire \bidir_PAD2CORE[42] ;
 wire \bidir_PAD2CORE[43] ;
 wire \bidir_PAD2CORE[44] ;
 wire \bidir_PAD2CORE[45] ;
 wire \bidir_PAD2CORE[46] ;
 wire \bidir_PAD2CORE[47] ;
 wire \bidir_PAD2CORE[48] ;
 wire \bidir_PAD2CORE[49] ;
 wire \bidir_PAD2CORE[4] ;
 wire \bidir_PAD2CORE[50] ;
 wire \bidir_PAD2CORE[51] ;
 wire \bidir_PAD2CORE[52] ;
 wire \bidir_PAD2CORE[53] ;
 wire \bidir_PAD2CORE[5] ;
 wire \bidir_PAD2CORE[6] ;
 wire \bidir_PAD2CORE[7] ;
 wire \bidir_PAD2CORE[8] ;
 wire \bidir_PAD2CORE[9] ;
 wire boot_rom_en;
 wire \bus_addr[0] ;
 wire \bus_addr[1] ;
 wire \bus_addr[2] ;
 wire \bus_addr[3] ;
 wire \bus_addr[4] ;
 wire \bus_addr[5] ;
 wire bus_cyc;
 wire \bus_data_gpios[0] ;
 wire \bus_data_gpios[1] ;
 wire \bus_data_gpios[2] ;
 wire \bus_data_gpios[3] ;
 wire \bus_data_gpios[4] ;
 wire \bus_data_gpios[5] ;
 wire \bus_data_gpios[6] ;
 wire \bus_data_gpios[7] ;
 wire \bus_data_out[0] ;
 wire \bus_data_out[1] ;
 wire \bus_data_out[2] ;
 wire \bus_data_out[3] ;
 wire \bus_data_out[4] ;
 wire \bus_data_out[5] ;
 wire \bus_data_out[6] ;
 wire \bus_data_out[7] ;
 wire \bus_data_serial_ports[0] ;
 wire \bus_data_serial_ports[1] ;
 wire \bus_data_serial_ports[2] ;
 wire \bus_data_serial_ports[3] ;
 wire \bus_data_serial_ports[4] ;
 wire \bus_data_serial_ports[5] ;
 wire \bus_data_serial_ports[6] ;
 wire \bus_data_serial_ports[7] ;
 wire \bus_data_sid[0] ;
 wire \bus_data_sid[1] ;
 wire \bus_data_sid[2] ;
 wire \bus_data_sid[3] ;
 wire \bus_data_sid[4] ;
 wire \bus_data_sid[5] ;
 wire \bus_data_sid[6] ;
 wire \bus_data_sid[7] ;
 wire \bus_data_timers[0] ;
 wire \bus_data_timers[1] ;
 wire \bus_data_timers[2] ;
 wire \bus_data_timers[3] ;
 wire \bus_data_timers[4] ;
 wire \bus_data_timers[5] ;
 wire \bus_data_timers[6] ;
 wire \bus_data_timers[7] ;
 wire bus_we_gpios;
 wire bus_we_serial_ports;
 wire bus_we_sid;
 wire bus_we_timers;
 wire clk_PAD2CORE;
 wire \const_zero[0] ;
 wire \const_zero[1] ;
 wire \const_zero[2] ;
 wire \const_zero[3] ;
 wire irq0;
 wire irq1;
 wire irq2;
 wire irq3;
 wire irq5;
 wire irq6;
 wire irq7;
 wire \last_addr[0] ;
 wire \last_addr[10] ;
 wire \last_addr[11] ;
 wire \last_addr[12] ;
 wire \last_addr[13] ;
 wire \last_addr[14] ;
 wire \last_addr[15] ;
 wire \last_addr[1] ;
 wire \last_addr[2] ;
 wire \last_addr[3] ;
 wire \last_addr[4] ;
 wire \last_addr[5] ;
 wire \last_addr[6] ;
 wire \last_addr[7] ;
 wire \last_addr[8] ;
 wire \last_addr[9] ;
 wire le_hi_act;
 wire le_lo_act;
 wire pwm0;
 wire pwm1;
 wire pwm2;
 wire \ram_bus_in[0] ;
 wire \ram_bus_in[1] ;
 wire \ram_bus_in[2] ;
 wire \ram_bus_in[3] ;
 wire \ram_bus_in[4] ;
 wire \ram_bus_in[5] ;
 wire \ram_bus_in[6] ;
 wire \ram_bus_in[7] ;
 wire ram_enabled;
 wire \requested_addr[0] ;
 wire \requested_addr[10] ;
 wire \requested_addr[11] ;
 wire \requested_addr[12] ;
 wire \requested_addr[13] ;
 wire \requested_addr[14] ;
 wire \requested_addr[15] ;
 wire \requested_addr[1] ;
 wire \requested_addr[2] ;
 wire \requested_addr[3] ;
 wire \requested_addr[4] ;
 wire \requested_addr[5] ;
 wire \requested_addr[6] ;
 wire \requested_addr[7] ;
 wire \requested_addr[8] ;
 wire \requested_addr[9] ;
 wire reset;
 wire \rom_bus_in[0] ;
 wire \rom_bus_in[1] ;
 wire \rom_bus_in[2] ;
 wire \rom_bus_in[3] ;
 wire \rom_bus_in[4] ;
 wire \rom_bus_in[5] ;
 wire \rom_bus_in[6] ;
 wire \rom_bus_in[7] ;
 wire \rom_bus_out[0] ;
 wire \rom_bus_out[1] ;
 wire \rom_bus_out[2] ;
 wire \rom_bus_out[3] ;
 wire \rom_bus_out[4] ;
 wire \rom_bus_out[5] ;
 wire \rom_bus_out[6] ;
 wire \rom_bus_out[7] ;
 wire rst_n_PAD2CORE;
 wire tmr0_clk;
 wire tmr0_o;
 wire tmr1_clk;
 wire tmr1_o;

 avali_logo avali_logo ();
 gf180mcu_fd_io__bi_24t \bidir[0].pad  (.A(\bidir_CORE2PAD[0] ),
    .CS(\bidir_CORE2PAD_CS[0] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[0] ),
    .OE(\bidir_CORE2PAD_OE[0] ),
    .PAD(bidir_PAD[0]),
    .PD(\bidir_CORE2PAD_PD[0] ),
    .PU(\bidir_CORE2PAD_PU[0] ),
    .SL(\bidir_CORE2PAD_SL[0] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[0] ));
 gf180mcu_fd_io__bi_24t \bidir[10].pad  (.A(\bidir_CORE2PAD[10] ),
    .CS(\bidir_CORE2PAD_CS[10] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[10] ),
    .OE(\bidir_CORE2PAD_OE[10] ),
    .PAD(bidir_PAD[10]),
    .PD(\bidir_CORE2PAD_PD[10] ),
    .PU(\bidir_CORE2PAD_PU[10] ),
    .SL(\bidir_CORE2PAD_SL[10] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[10] ));
 gf180mcu_fd_io__bi_24t \bidir[11].pad  (.A(\bidir_CORE2PAD[11] ),
    .CS(\bidir_CORE2PAD_CS[11] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[11] ),
    .OE(\bidir_CORE2PAD_OE[11] ),
    .PAD(bidir_PAD[11]),
    .PD(\bidir_CORE2PAD_PD[11] ),
    .PU(\bidir_CORE2PAD_PU[11] ),
    .SL(\bidir_CORE2PAD_SL[11] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[11] ));
 gf180mcu_fd_io__bi_24t \bidir[12].pad  (.A(\bidir_CORE2PAD[12] ),
    .CS(\bidir_CORE2PAD_CS[12] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[12] ),
    .OE(\bidir_CORE2PAD_OE[12] ),
    .PAD(bidir_PAD[12]),
    .PD(\bidir_CORE2PAD_PD[12] ),
    .PU(\bidir_CORE2PAD_PU[12] ),
    .SL(\bidir_CORE2PAD_SL[12] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[12] ));
 gf180mcu_fd_io__bi_24t \bidir[13].pad  (.A(\bidir_CORE2PAD[13] ),
    .CS(\bidir_CORE2PAD_CS[13] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[13] ),
    .OE(\bidir_CORE2PAD_OE[13] ),
    .PAD(bidir_PAD[13]),
    .PD(\bidir_CORE2PAD_PD[13] ),
    .PU(\bidir_CORE2PAD_PU[13] ),
    .SL(\bidir_CORE2PAD_SL[13] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[13] ));
 gf180mcu_fd_io__bi_24t \bidir[14].pad  (.A(\bidir_CORE2PAD[14] ),
    .CS(\bidir_CORE2PAD_CS[14] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[14] ),
    .OE(\bidir_CORE2PAD_OE[14] ),
    .PAD(bidir_PAD[14]),
    .PD(\bidir_CORE2PAD_PD[14] ),
    .PU(\bidir_CORE2PAD_PU[14] ),
    .SL(\bidir_CORE2PAD_SL[14] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[14] ));
 gf180mcu_fd_io__bi_24t \bidir[15].pad  (.A(\bidir_CORE2PAD[15] ),
    .CS(\bidir_CORE2PAD_CS[15] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[15] ),
    .OE(\bidir_CORE2PAD_OE[15] ),
    .PAD(bidir_PAD[15]),
    .PD(\bidir_CORE2PAD_PD[15] ),
    .PU(\bidir_CORE2PAD_PU[15] ),
    .SL(\bidir_CORE2PAD_SL[15] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[15] ));
 gf180mcu_fd_io__bi_24t \bidir[16].pad  (.A(\bidir_CORE2PAD[16] ),
    .CS(\bidir_CORE2PAD_CS[16] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[16] ),
    .OE(\bidir_CORE2PAD_OE[16] ),
    .PAD(bidir_PAD[16]),
    .PD(\bidir_CORE2PAD_PD[16] ),
    .PU(\bidir_CORE2PAD_PU[16] ),
    .SL(\bidir_CORE2PAD_SL[16] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[16] ));
 gf180mcu_fd_io__bi_24t \bidir[17].pad  (.A(\bidir_CORE2PAD[17] ),
    .CS(\bidir_CORE2PAD_CS[17] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[17] ),
    .OE(\bidir_CORE2PAD_OE[17] ),
    .PAD(bidir_PAD[17]),
    .PD(\bidir_CORE2PAD_PD[17] ),
    .PU(\bidir_CORE2PAD_PU[17] ),
    .SL(\bidir_CORE2PAD_SL[17] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[17] ));
 gf180mcu_fd_io__bi_24t \bidir[18].pad  (.A(\bidir_CORE2PAD[18] ),
    .CS(\bidir_CORE2PAD_CS[18] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[18] ),
    .OE(\bidir_CORE2PAD_OE[18] ),
    .PAD(bidir_PAD[18]),
    .PD(\bidir_CORE2PAD_PD[18] ),
    .PU(\bidir_CORE2PAD_PU[18] ),
    .SL(\bidir_CORE2PAD_SL[18] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[18] ));
 gf180mcu_fd_io__bi_24t \bidir[19].pad  (.A(\bidir_CORE2PAD[19] ),
    .CS(\bidir_CORE2PAD_CS[19] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[19] ),
    .OE(\bidir_CORE2PAD_OE[19] ),
    .PAD(bidir_PAD[19]),
    .PD(\bidir_CORE2PAD_PD[19] ),
    .PU(\bidir_CORE2PAD_PU[19] ),
    .SL(\bidir_CORE2PAD_SL[19] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[19] ));
 gf180mcu_fd_io__bi_24t \bidir[1].pad  (.A(\bidir_CORE2PAD[1] ),
    .CS(\bidir_CORE2PAD_CS[1] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[1] ),
    .OE(\bidir_CORE2PAD_OE[1] ),
    .PAD(bidir_PAD[1]),
    .PD(\bidir_CORE2PAD_PD[1] ),
    .PU(\bidir_CORE2PAD_PU[1] ),
    .SL(\bidir_CORE2PAD_SL[1] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[1] ));
 gf180mcu_fd_io__bi_24t \bidir[20].pad  (.A(\bidir_CORE2PAD[20] ),
    .CS(\bidir_CORE2PAD_CS[20] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[20] ),
    .OE(\bidir_CORE2PAD_OE[20] ),
    .PAD(bidir_PAD[20]),
    .PD(\bidir_CORE2PAD_PD[20] ),
    .PU(\bidir_CORE2PAD_PU[20] ),
    .SL(\bidir_CORE2PAD_SL[20] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[20] ));
 gf180mcu_fd_io__bi_24t \bidir[21].pad  (.A(\bidir_CORE2PAD[21] ),
    .CS(\bidir_CORE2PAD_CS[21] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[21] ),
    .OE(\bidir_CORE2PAD_OE[21] ),
    .PAD(bidir_PAD[21]),
    .PD(\bidir_CORE2PAD_PD[21] ),
    .PU(\bidir_CORE2PAD_PU[21] ),
    .SL(\bidir_CORE2PAD_SL[21] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[21] ));
 gf180mcu_fd_io__bi_24t \bidir[22].pad  (.A(\bidir_CORE2PAD[22] ),
    .CS(\bidir_CORE2PAD_CS[22] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[22] ),
    .OE(\bidir_CORE2PAD_OE[22] ),
    .PAD(bidir_PAD[22]),
    .PD(\bidir_CORE2PAD_PD[22] ),
    .PU(\bidir_CORE2PAD_PU[22] ),
    .SL(\bidir_CORE2PAD_SL[22] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[22] ));
 gf180mcu_fd_io__bi_24t \bidir[23].pad  (.A(\bidir_CORE2PAD[23] ),
    .CS(\bidir_CORE2PAD_CS[23] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[23] ),
    .OE(\bidir_CORE2PAD_OE[23] ),
    .PAD(bidir_PAD[23]),
    .PD(\bidir_CORE2PAD_PD[23] ),
    .PU(\bidir_CORE2PAD_PU[23] ),
    .SL(\bidir_CORE2PAD_SL[23] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[23] ));
 gf180mcu_fd_io__bi_24t \bidir[24].pad  (.A(\bidir_CORE2PAD[24] ),
    .CS(\bidir_CORE2PAD_CS[24] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[24] ),
    .OE(\bidir_CORE2PAD_OE[24] ),
    .PAD(bidir_PAD[24]),
    .PD(\bidir_CORE2PAD_PD[24] ),
    .PU(\bidir_CORE2PAD_PU[24] ),
    .SL(\bidir_CORE2PAD_SL[24] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[24] ));
 gf180mcu_fd_io__bi_24t \bidir[25].pad  (.A(\bidir_CORE2PAD[25] ),
    .CS(\bidir_CORE2PAD_CS[25] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[25] ),
    .OE(\bidir_CORE2PAD_OE[25] ),
    .PAD(bidir_PAD[25]),
    .PD(\bidir_CORE2PAD_PD[25] ),
    .PU(\bidir_CORE2PAD_PU[25] ),
    .SL(\bidir_CORE2PAD_SL[25] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[25] ));
 gf180mcu_fd_io__bi_24t \bidir[26].pad  (.A(\bidir_CORE2PAD[26] ),
    .CS(\bidir_CORE2PAD_CS[26] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[26] ),
    .OE(\bidir_CORE2PAD_OE[26] ),
    .PAD(bidir_PAD[26]),
    .PD(\bidir_CORE2PAD_PD[26] ),
    .PU(\bidir_CORE2PAD_PU[26] ),
    .SL(\bidir_CORE2PAD_SL[26] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[26] ));
 gf180mcu_fd_io__bi_24t \bidir[27].pad  (.A(\bidir_CORE2PAD[27] ),
    .CS(\bidir_CORE2PAD_CS[27] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[27] ),
    .OE(\bidir_CORE2PAD_OE[27] ),
    .PAD(bidir_PAD[27]),
    .PD(\bidir_CORE2PAD_PD[27] ),
    .PU(\bidir_CORE2PAD_PU[27] ),
    .SL(\bidir_CORE2PAD_SL[27] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[27] ));
 gf180mcu_fd_io__bi_24t \bidir[28].pad  (.A(\bidir_CORE2PAD[28] ),
    .CS(\bidir_CORE2PAD_CS[28] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[28] ),
    .OE(\bidir_CORE2PAD_OE[28] ),
    .PAD(bidir_PAD[28]),
    .PD(\bidir_CORE2PAD_PD[28] ),
    .PU(\bidir_CORE2PAD_PU[28] ),
    .SL(\bidir_CORE2PAD_SL[28] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[28] ));
 gf180mcu_fd_io__bi_24t \bidir[29].pad  (.A(\bidir_CORE2PAD[29] ),
    .CS(\bidir_CORE2PAD_CS[29] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[29] ),
    .OE(\bidir_CORE2PAD_OE[29] ),
    .PAD(bidir_PAD[29]),
    .PD(\bidir_CORE2PAD_PD[29] ),
    .PU(\bidir_CORE2PAD_PU[29] ),
    .SL(\bidir_CORE2PAD_SL[29] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[29] ));
 gf180mcu_fd_io__bi_24t \bidir[2].pad  (.A(\bidir_CORE2PAD[2] ),
    .CS(\bidir_CORE2PAD_CS[2] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[2] ),
    .OE(\bidir_CORE2PAD_OE[2] ),
    .PAD(bidir_PAD[2]),
    .PD(\bidir_CORE2PAD_PD[2] ),
    .PU(\bidir_CORE2PAD_PU[2] ),
    .SL(\bidir_CORE2PAD_SL[2] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[2] ));
 gf180mcu_fd_io__bi_24t \bidir[30].pad  (.A(\bidir_CORE2PAD[30] ),
    .CS(\bidir_CORE2PAD_CS[30] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[30] ),
    .OE(\bidir_CORE2PAD_OE[30] ),
    .PAD(bidir_PAD[30]),
    .PD(\bidir_CORE2PAD_PD[30] ),
    .PU(\bidir_CORE2PAD_PU[30] ),
    .SL(\bidir_CORE2PAD_SL[30] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[30] ));
 gf180mcu_fd_io__bi_24t \bidir[31].pad  (.A(\bidir_CORE2PAD[31] ),
    .CS(\bidir_CORE2PAD_CS[31] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[31] ),
    .OE(\bidir_CORE2PAD_OE[31] ),
    .PAD(bidir_PAD[31]),
    .PD(\bidir_CORE2PAD_PD[31] ),
    .PU(\bidir_CORE2PAD_PU[31] ),
    .SL(\bidir_CORE2PAD_SL[31] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[31] ));
 gf180mcu_fd_io__bi_24t \bidir[32].pad  (.A(\bidir_CORE2PAD[32] ),
    .CS(\bidir_CORE2PAD_CS[32] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[32] ),
    .OE(\bidir_CORE2PAD_OE[32] ),
    .PAD(bidir_PAD[32]),
    .PD(\bidir_CORE2PAD_PD[32] ),
    .PU(\bidir_CORE2PAD_PU[32] ),
    .SL(\bidir_CORE2PAD_SL[32] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[32] ));
 gf180mcu_fd_io__bi_24t \bidir[33].pad  (.A(\bidir_CORE2PAD[33] ),
    .CS(\bidir_CORE2PAD_CS[33] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[33] ),
    .OE(\bidir_CORE2PAD_OE[33] ),
    .PAD(bidir_PAD[33]),
    .PD(\bidir_CORE2PAD_PD[33] ),
    .PU(\bidir_CORE2PAD_PU[33] ),
    .SL(\bidir_CORE2PAD_SL[33] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[33] ));
 gf180mcu_fd_io__bi_24t \bidir[34].pad  (.A(\bidir_CORE2PAD[34] ),
    .CS(\bidir_CORE2PAD_CS[34] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[34] ),
    .OE(\bidir_CORE2PAD_OE[34] ),
    .PAD(bidir_PAD[34]),
    .PD(\bidir_CORE2PAD_PD[34] ),
    .PU(\bidir_CORE2PAD_PU[34] ),
    .SL(\bidir_CORE2PAD_SL[34] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[34] ));
 gf180mcu_fd_io__bi_24t \bidir[35].pad  (.A(\bidir_CORE2PAD[35] ),
    .CS(\bidir_CORE2PAD_CS[35] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[35] ),
    .OE(\bidir_CORE2PAD_OE[35] ),
    .PAD(bidir_PAD[35]),
    .PD(\bidir_CORE2PAD_PD[35] ),
    .PU(\bidir_CORE2PAD_PU[35] ),
    .SL(\bidir_CORE2PAD_SL[35] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[35] ));
 gf180mcu_fd_io__bi_24t \bidir[36].pad  (.A(\bidir_CORE2PAD[36] ),
    .CS(\bidir_CORE2PAD_CS[36] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[36] ),
    .OE(\bidir_CORE2PAD_OE[36] ),
    .PAD(bidir_PAD[36]),
    .PD(\bidir_CORE2PAD_PD[36] ),
    .PU(\bidir_CORE2PAD_PU[36] ),
    .SL(\bidir_CORE2PAD_SL[36] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[36] ));
 gf180mcu_fd_io__bi_24t \bidir[37].pad  (.A(\bidir_CORE2PAD[37] ),
    .CS(\bidir_CORE2PAD_CS[37] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[37] ),
    .OE(\bidir_CORE2PAD_OE[37] ),
    .PAD(bidir_PAD[37]),
    .PD(\bidir_CORE2PAD_PD[37] ),
    .PU(\bidir_CORE2PAD_PU[37] ),
    .SL(\bidir_CORE2PAD_SL[37] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[37] ));
 gf180mcu_fd_io__bi_24t \bidir[38].pad  (.A(\bidir_CORE2PAD[38] ),
    .CS(\bidir_CORE2PAD_CS[38] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[38] ),
    .OE(\bidir_CORE2PAD_OE[38] ),
    .PAD(bidir_PAD[38]),
    .PD(\bidir_CORE2PAD_PD[38] ),
    .PU(\bidir_CORE2PAD_PU[38] ),
    .SL(\bidir_CORE2PAD_SL[38] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[38] ));
 gf180mcu_fd_io__bi_24t \bidir[39].pad  (.A(\bidir_CORE2PAD[39] ),
    .CS(\bidir_CORE2PAD_CS[39] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[39] ),
    .OE(\bidir_CORE2PAD_OE[39] ),
    .PAD(bidir_PAD[39]),
    .PD(\bidir_CORE2PAD_PD[39] ),
    .PU(\bidir_CORE2PAD_PU[39] ),
    .SL(\bidir_CORE2PAD_SL[39] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[39] ));
 gf180mcu_fd_io__bi_24t \bidir[3].pad  (.A(\bidir_CORE2PAD[3] ),
    .CS(\bidir_CORE2PAD_CS[3] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[3] ),
    .OE(\bidir_CORE2PAD_OE[3] ),
    .PAD(bidir_PAD[3]),
    .PD(\bidir_CORE2PAD_PD[3] ),
    .PU(\bidir_CORE2PAD_PU[3] ),
    .SL(\bidir_CORE2PAD_SL[3] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[3] ));
 gf180mcu_fd_io__bi_24t \bidir[40].pad  (.A(\bidir_CORE2PAD[40] ),
    .CS(\bidir_CORE2PAD_CS[40] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[40] ),
    .OE(\bidir_CORE2PAD_OE[40] ),
    .PAD(bidir_PAD[40]),
    .PD(\bidir_CORE2PAD_PD[40] ),
    .PU(\bidir_CORE2PAD_PU[40] ),
    .SL(\bidir_CORE2PAD_SL[40] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[40] ));
 gf180mcu_fd_io__bi_24t \bidir[41].pad  (.A(\bidir_CORE2PAD[41] ),
    .CS(\bidir_CORE2PAD_CS[41] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[41] ),
    .OE(\bidir_CORE2PAD_OE[41] ),
    .PAD(bidir_PAD[41]),
    .PD(\bidir_CORE2PAD_PD[41] ),
    .PU(\bidir_CORE2PAD_PU[41] ),
    .SL(\bidir_CORE2PAD_SL[41] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[41] ));
 gf180mcu_fd_io__bi_24t \bidir[42].pad  (.A(\bidir_CORE2PAD[42] ),
    .CS(\bidir_CORE2PAD_CS[42] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[42] ),
    .OE(\bidir_CORE2PAD_OE[42] ),
    .PAD(bidir_PAD[42]),
    .PD(\bidir_CORE2PAD_PD[42] ),
    .PU(\bidir_CORE2PAD_PU[42] ),
    .SL(\bidir_CORE2PAD_SL[42] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[42] ));
 gf180mcu_fd_io__bi_24t \bidir[43].pad  (.A(\bidir_CORE2PAD[43] ),
    .CS(\bidir_CORE2PAD_CS[43] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[43] ),
    .OE(\bidir_CORE2PAD_OE[43] ),
    .PAD(bidir_PAD[43]),
    .PD(\bidir_CORE2PAD_PD[43] ),
    .PU(\bidir_CORE2PAD_PU[43] ),
    .SL(\bidir_CORE2PAD_SL[43] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[43] ));
 gf180mcu_fd_io__bi_24t \bidir[44].pad  (.A(\bidir_CORE2PAD[44] ),
    .CS(\bidir_CORE2PAD_CS[44] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[44] ),
    .OE(\bidir_CORE2PAD_OE[44] ),
    .PAD(bidir_PAD[44]),
    .PD(\bidir_CORE2PAD_PD[44] ),
    .PU(\bidir_CORE2PAD_PU[44] ),
    .SL(\bidir_CORE2PAD_SL[44] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[44] ));
 gf180mcu_fd_io__bi_24t \bidir[45].pad  (.A(\bidir_CORE2PAD[45] ),
    .CS(\bidir_CORE2PAD_CS[45] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[45] ),
    .OE(\bidir_CORE2PAD_OE[45] ),
    .PAD(bidir_PAD[45]),
    .PD(\bidir_CORE2PAD_PD[45] ),
    .PU(\bidir_CORE2PAD_PU[45] ),
    .SL(\bidir_CORE2PAD_SL[45] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[45] ));
 gf180mcu_fd_io__bi_24t \bidir[46].pad  (.A(\bidir_CORE2PAD[46] ),
    .CS(\bidir_CORE2PAD_CS[46] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[46] ),
    .OE(\bidir_CORE2PAD_OE[46] ),
    .PAD(bidir_PAD[46]),
    .PD(\bidir_CORE2PAD_PD[46] ),
    .PU(\bidir_CORE2PAD_PU[46] ),
    .SL(\bidir_CORE2PAD_SL[46] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[46] ));
 gf180mcu_fd_io__bi_24t \bidir[47].pad  (.A(\bidir_CORE2PAD[47] ),
    .CS(\bidir_CORE2PAD_CS[47] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[47] ),
    .OE(\bidir_CORE2PAD_OE[47] ),
    .PAD(bidir_PAD[47]),
    .PD(\bidir_CORE2PAD_PD[47] ),
    .PU(\bidir_CORE2PAD_PU[47] ),
    .SL(\bidir_CORE2PAD_SL[47] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[47] ));
 gf180mcu_fd_io__bi_24t \bidir[48].pad  (.A(\bidir_CORE2PAD[48] ),
    .CS(\bidir_CORE2PAD_CS[48] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[48] ),
    .OE(\bidir_CORE2PAD_OE[48] ),
    .PAD(bidir_PAD[48]),
    .PD(\bidir_CORE2PAD_PD[48] ),
    .PU(\bidir_CORE2PAD_PU[48] ),
    .SL(\bidir_CORE2PAD_SL[48] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[48] ));
 gf180mcu_fd_io__bi_24t \bidir[49].pad  (.A(\bidir_CORE2PAD[49] ),
    .CS(\bidir_CORE2PAD_CS[49] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[49] ),
    .OE(\bidir_CORE2PAD_OE[49] ),
    .PAD(bidir_PAD[49]),
    .PD(\bidir_CORE2PAD_PD[49] ),
    .PU(\bidir_CORE2PAD_PU[49] ),
    .SL(\bidir_CORE2PAD_SL[49] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[49] ));
 gf180mcu_fd_io__bi_24t \bidir[4].pad  (.A(\bidir_CORE2PAD[4] ),
    .CS(\bidir_CORE2PAD_CS[4] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[4] ),
    .OE(\bidir_CORE2PAD_OE[4] ),
    .PAD(bidir_PAD[4]),
    .PD(\bidir_CORE2PAD_PD[4] ),
    .PU(\bidir_CORE2PAD_PU[4] ),
    .SL(\bidir_CORE2PAD_SL[4] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[4] ));
 gf180mcu_fd_io__bi_24t \bidir[50].pad  (.A(\bidir_CORE2PAD[50] ),
    .CS(\bidir_CORE2PAD_CS[50] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[50] ),
    .OE(\bidir_CORE2PAD_OE[50] ),
    .PAD(bidir_PAD[50]),
    .PD(\bidir_CORE2PAD_PD[50] ),
    .PU(\bidir_CORE2PAD_PU[50] ),
    .SL(\bidir_CORE2PAD_SL[50] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[50] ));
 gf180mcu_fd_io__bi_24t \bidir[51].pad  (.A(\bidir_CORE2PAD[51] ),
    .CS(\bidir_CORE2PAD_CS[51] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[51] ),
    .OE(\bidir_CORE2PAD_OE[51] ),
    .PAD(bidir_PAD[51]),
    .PD(\bidir_CORE2PAD_PD[51] ),
    .PU(\bidir_CORE2PAD_PU[51] ),
    .SL(\bidir_CORE2PAD_SL[51] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[51] ));
 gf180mcu_fd_io__bi_24t \bidir[52].pad  (.A(\bidir_CORE2PAD[52] ),
    .CS(\bidir_CORE2PAD_CS[52] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[52] ),
    .OE(\bidir_CORE2PAD_OE[52] ),
    .PAD(bidir_PAD[52]),
    .PD(\bidir_CORE2PAD_PD[52] ),
    .PU(\bidir_CORE2PAD_PU[52] ),
    .SL(\bidir_CORE2PAD_SL[52] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[52] ));
 gf180mcu_fd_io__bi_24t \bidir[53].pad  (.A(\bidir_CORE2PAD[53] ),
    .CS(\bidir_CORE2PAD_CS[53] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[53] ),
    .OE(\bidir_CORE2PAD_OE[53] ),
    .PAD(bidir_PAD[53]),
    .PD(\bidir_CORE2PAD_PD[53] ),
    .PU(\bidir_CORE2PAD_PU[53] ),
    .SL(\bidir_CORE2PAD_SL[53] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[53] ));
 gf180mcu_fd_io__bi_24t \bidir[5].pad  (.A(\bidir_CORE2PAD[5] ),
    .CS(\bidir_CORE2PAD_CS[5] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[5] ),
    .OE(\bidir_CORE2PAD_OE[5] ),
    .PAD(bidir_PAD[5]),
    .PD(\bidir_CORE2PAD_PD[5] ),
    .PU(\bidir_CORE2PAD_PU[5] ),
    .SL(\bidir_CORE2PAD_SL[5] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[5] ));
 gf180mcu_fd_io__bi_24t \bidir[6].pad  (.A(\bidir_CORE2PAD[6] ),
    .CS(\bidir_CORE2PAD_CS[6] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[6] ),
    .OE(\bidir_CORE2PAD_OE[6] ),
    .PAD(bidir_PAD[6]),
    .PD(\bidir_CORE2PAD_PD[6] ),
    .PU(\bidir_CORE2PAD_PU[6] ),
    .SL(\bidir_CORE2PAD_SL[6] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[6] ));
 gf180mcu_fd_io__bi_24t \bidir[7].pad  (.A(\bidir_CORE2PAD[7] ),
    .CS(\bidir_CORE2PAD_CS[7] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[7] ),
    .OE(\bidir_CORE2PAD_OE[7] ),
    .PAD(bidir_PAD[7]),
    .PD(\bidir_CORE2PAD_PD[7] ),
    .PU(\bidir_CORE2PAD_PU[7] ),
    .SL(\bidir_CORE2PAD_SL[7] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[7] ));
 gf180mcu_fd_io__bi_24t \bidir[8].pad  (.A(\bidir_CORE2PAD[8] ),
    .CS(\bidir_CORE2PAD_CS[8] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[8] ),
    .OE(\bidir_CORE2PAD_OE[8] ),
    .PAD(bidir_PAD[8]),
    .PD(\bidir_CORE2PAD_PD[8] ),
    .PU(\bidir_CORE2PAD_PU[8] ),
    .SL(\bidir_CORE2PAD_SL[8] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[8] ));
 gf180mcu_fd_io__bi_24t \bidir[9].pad  (.A(\bidir_CORE2PAD[9] ),
    .CS(\bidir_CORE2PAD_CS[9] ),
    .DVDD(VDD),
    .DVSS(VSS),
    .IE(\bidir_CORE2PAD_IE[9] ),
    .OE(\bidir_CORE2PAD_OE[9] ),
    .PAD(bidir_PAD[9]),
    .PD(\bidir_CORE2PAD_PD[9] ),
    .PU(\bidir_CORE2PAD_PU[9] ),
    .SL(\bidir_CORE2PAD_SL[9] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(\bidir_PAD2CORE[9] ));
 boot_rom boot_rom (.VDD(VDD),
    .VSS(VSS),
    .clk_i(clk_PAD2CORE),
    .rst(reset),
    .bus_out({\rom_bus_in[7] ,
    \rom_bus_in[6] ,
    \rom_bus_in[5] ,
    \rom_bus_in[4] ,
    \rom_bus_in[3] ,
    \rom_bus_in[2] ,
    \rom_bus_in[1] ,
    \rom_bus_in[0] }),
    .last_addr({\last_addr[7] ,
    \last_addr[6] ,
    \last_addr[5] ,
    \last_addr[4] ,
    \last_addr[3] ,
    \last_addr[2] ,
    \last_addr[1] ,
    \last_addr[0] }));
 gf180mcu_ws_ip__id chip_id ();
 gf180mcu_fd_io__in_s clk_pad (.DVDD(VDD),
    .DVSS(VSS),
    .PAD(clk_PAD),
    .PD(\const_zero[3] ),
    .PU(\const_zero[2] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(clk_PAD2CORE));
 gf180mcu_ws_io__dvdd dvdd_east_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VSS(VSS));
 gf180mcu_ws_io__dvdd dvdd_east_1 (.DVDD(VDD),
    .DVSS(VSS),
    .VSS(VSS));
 gf180mcu_ws_io__dvdd dvdd_east_2 (.DVDD(VDD),
    .DVSS(VSS),
    .VSS(VSS));
 gf180mcu_ws_io__dvdd dvdd_east_3 (.DVDD(VDD),
    .DVSS(VSS),
    .VSS(VSS));
 gf180mcu_ws_io__dvdd dvdd_west_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VSS(VSS));
 gf180mcu_ws_io__dvdd dvdd_west_1 (.DVDD(VDD),
    .DVSS(VSS),
    .VSS(VSS));
 gf180mcu_ws_io__dvdd dvdd_west_2 (.DVDD(VDD),
    .DVSS(VSS),
    .VSS(VSS));
 gf180mcu_ws_io__dvdd dvdd_west_3 (.DVDD(VDD),
    .DVSS(VSS),
    .VSS(VSS));
 gf180mcu_ws_io__dvss dvss_east_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_ws_io__dvss dvss_east_1 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_ws_io__dvss dvss_east_2 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_ws_io__dvss dvss_east_3 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_fd_io__dvss dvss_north_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_fd_io__dvss dvss_south_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_ws_io__dvss dvss_west_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_ws_io__dvss dvss_west_1 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_ws_io__dvss dvss_west_2 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gf180mcu_ws_io__dvss dvss_west_3 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD));
 gpios gpios (.DAC_clk(DAC_clk),
    .DAC_d1(DAC_d1),
    .DAC_d2(DAC_d2),
    .DAC_le(DAC_le),
    .RXD(RXD),
    .TXD(TXD),
    .VDD(VDD),
    .VSS(VSS),
    .bus_cyc(bus_cyc),
    .bus_we(bus_we_gpios),
    .clk_i(clk_PAD2CORE),
    .irq0(irq0),
    .irq6(irq6),
    .irq7(irq7),
    .pwm0(pwm0),
    .pwm1(pwm1),
    .pwm2(pwm2),
    .rst(reset),
    .tmr0_clk(tmr0_clk),
    .tmr0_o(tmr0_o),
    .tmr1_clk(tmr1_clk),
    .tmr1_o(tmr1_o),
    .addr({\bus_addr[3] ,
    \bus_addr[2] ,
    \bus_addr[1] ,
    \bus_addr[0] }),
    .data_in({\bus_data_out[7] ,
    \bus_data_out[6] ,
    \bus_data_out[5] ,
    \bus_data_out[4] ,
    \bus_data_out[3] ,
    \bus_data_out[2] ,
    \bus_data_out[1] ,
    \bus_data_out[0] }),
    .data_out({\bus_data_gpios[7] ,
    \bus_data_gpios[6] ,
    \bus_data_gpios[5] ,
    \bus_data_gpios[4] ,
    \bus_data_gpios[3] ,
    \bus_data_gpios[2] ,
    \bus_data_gpios[1] ,
    \bus_data_gpios[0] }),
    .io_cs({\bidir_CORE2PAD_CS[34] ,
    \bidir_CORE2PAD_CS[33] ,
    \bidir_CORE2PAD_CS[32] ,
    \bidir_CORE2PAD_CS[31] ,
    \bidir_CORE2PAD_CS[30] ,
    \bidir_CORE2PAD_CS[29] ,
    \bidir_CORE2PAD_CS[28] ,
    \bidir_CORE2PAD_CS[27] ,
    \bidir_CORE2PAD_CS[26] ,
    \bidir_CORE2PAD_CS[25] ,
    \bidir_CORE2PAD_CS[24] ,
    \bidir_CORE2PAD_CS[23] ,
    \bidir_CORE2PAD_CS[22] ,
    \bidir_CORE2PAD_CS[21] ,
    \bidir_CORE2PAD_CS[20] ,
    \bidir_CORE2PAD_CS[19] }),
    .io_ie({\bidir_CORE2PAD_IE[34] ,
    \bidir_CORE2PAD_IE[33] ,
    \bidir_CORE2PAD_IE[32] ,
    \bidir_CORE2PAD_IE[31] ,
    \bidir_CORE2PAD_IE[30] ,
    \bidir_CORE2PAD_IE[29] ,
    \bidir_CORE2PAD_IE[28] ,
    \bidir_CORE2PAD_IE[27] ,
    \bidir_CORE2PAD_IE[26] ,
    \bidir_CORE2PAD_IE[25] ,
    \bidir_CORE2PAD_IE[24] ,
    \bidir_CORE2PAD_IE[23] ,
    \bidir_CORE2PAD_IE[22] ,
    \bidir_CORE2PAD_IE[21] ,
    \bidir_CORE2PAD_IE[20] ,
    \bidir_CORE2PAD_IE[19] }),
    .io_in({\bidir_PAD2CORE[34] ,
    \bidir_PAD2CORE[33] ,
    \bidir_PAD2CORE[32] ,
    \bidir_PAD2CORE[31] ,
    \bidir_PAD2CORE[30] ,
    \bidir_PAD2CORE[29] ,
    \bidir_PAD2CORE[28] ,
    \bidir_PAD2CORE[27] ,
    \bidir_PAD2CORE[26] ,
    \bidir_PAD2CORE[25] ,
    \bidir_PAD2CORE[24] ,
    \bidir_PAD2CORE[23] ,
    \bidir_PAD2CORE[22] ,
    \bidir_PAD2CORE[21] ,
    \bidir_PAD2CORE[20] ,
    \bidir_PAD2CORE[19] }),
    .io_oe({\bidir_CORE2PAD_OE[34] ,
    \bidir_CORE2PAD_OE[33] ,
    \bidir_CORE2PAD_OE[32] ,
    \bidir_CORE2PAD_OE[31] ,
    \bidir_CORE2PAD_OE[30] ,
    \bidir_CORE2PAD_OE[29] ,
    \bidir_CORE2PAD_OE[28] ,
    \bidir_CORE2PAD_OE[27] ,
    \bidir_CORE2PAD_OE[26] ,
    \bidir_CORE2PAD_OE[25] ,
    \bidir_CORE2PAD_OE[24] ,
    \bidir_CORE2PAD_OE[23] ,
    \bidir_CORE2PAD_OE[22] ,
    \bidir_CORE2PAD_OE[21] ,
    \bidir_CORE2PAD_OE[20] ,
    \bidir_CORE2PAD_OE[19] }),
    .io_out({\bidir_CORE2PAD[34] ,
    \bidir_CORE2PAD[33] ,
    \bidir_CORE2PAD[32] ,
    \bidir_CORE2PAD[31] ,
    \bidir_CORE2PAD[30] ,
    \bidir_CORE2PAD[29] ,
    \bidir_CORE2PAD[28] ,
    \bidir_CORE2PAD[27] ,
    \bidir_CORE2PAD[26] ,
    \bidir_CORE2PAD[25] ,
    \bidir_CORE2PAD[24] ,
    \bidir_CORE2PAD[23] ,
    \bidir_CORE2PAD[22] ,
    \bidir_CORE2PAD[21] ,
    \bidir_CORE2PAD[20] ,
    \bidir_CORE2PAD[19] }),
    .io_pd({\bidir_CORE2PAD_PD[34] ,
    \bidir_CORE2PAD_PD[33] ,
    \bidir_CORE2PAD_PD[32] ,
    \bidir_CORE2PAD_PD[31] ,
    \bidir_CORE2PAD_PD[30] ,
    \bidir_CORE2PAD_PD[29] ,
    \bidir_CORE2PAD_PD[28] ,
    \bidir_CORE2PAD_PD[27] ,
    \bidir_CORE2PAD_PD[26] ,
    \bidir_CORE2PAD_PD[25] ,
    \bidir_CORE2PAD_PD[24] ,
    \bidir_CORE2PAD_PD[23] ,
    \bidir_CORE2PAD_PD[22] ,
    \bidir_CORE2PAD_PD[21] ,
    \bidir_CORE2PAD_PD[20] ,
    \bidir_CORE2PAD_PD[19] }),
    .io_pu({\bidir_CORE2PAD_PU[34] ,
    \bidir_CORE2PAD_PU[33] ,
    \bidir_CORE2PAD_PU[32] ,
    \bidir_CORE2PAD_PU[31] ,
    \bidir_CORE2PAD_PU[30] ,
    \bidir_CORE2PAD_PU[29] ,
    \bidir_CORE2PAD_PU[28] ,
    \bidir_CORE2PAD_PU[27] ,
    \bidir_CORE2PAD_PU[26] ,
    \bidir_CORE2PAD_PU[25] ,
    \bidir_CORE2PAD_PU[24] ,
    \bidir_CORE2PAD_PU[23] ,
    \bidir_CORE2PAD_PU[22] ,
    \bidir_CORE2PAD_PU[21] ,
    \bidir_CORE2PAD_PU[20] ,
    \bidir_CORE2PAD_PU[19] }),
    .io_sl({\bidir_CORE2PAD_SL[34] ,
    \bidir_CORE2PAD_SL[33] ,
    \bidir_CORE2PAD_SL[32] ,
    \bidir_CORE2PAD_SL[31] ,
    \bidir_CORE2PAD_SL[30] ,
    \bidir_CORE2PAD_SL[29] ,
    \bidir_CORE2PAD_SL[28] ,
    \bidir_CORE2PAD_SL[27] ,
    \bidir_CORE2PAD_SL[26] ,
    \bidir_CORE2PAD_SL[25] ,
    \bidir_CORE2PAD_SL[24] ,
    \bidir_CORE2PAD_SL[23] ,
    \bidir_CORE2PAD_SL[22] ,
    \bidir_CORE2PAD_SL[21] ,
    \bidir_CORE2PAD_SL[20] ,
    \bidir_CORE2PAD_SL[19] }));
 ram_controller ram_controller (.CEN_all(CEN_all),
    .GWEN_0(GWEN_0),
    .GWEN_1(GWEN_1),
    .GWEN_2(GWEN_2),
    .GWEN_3(GWEN_3),
    .GWEN_4(GWEN_4),
    .GWEN_5(GWEN_5),
    .GWEN_6(GWEN_6),
    .GWEN_7(GWEN_7),
    .VDD(VDD),
    .VSS(VSS),
    .WEb_ram(WEb_ram),
    .clk_i(clk_PAD2CORE),
    .ram_enabled(ram_enabled),
    .rst(reset),
    .A_all({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D_all({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q0({\Q0[7] ,
    \Q0[6] ,
    \Q0[5] ,
    \Q0[4] ,
    \Q0[3] ,
    \Q0[2] ,
    \Q0[1] ,
    \Q0[0] }),
    .Q1({\Q1[7] ,
    \Q1[6] ,
    \Q1[5] ,
    \Q1[4] ,
    \Q1[3] ,
    \Q1[2] ,
    \Q1[1] ,
    \Q1[0] }),
    .Q2({\Q2[7] ,
    \Q2[6] ,
    \Q2[5] ,
    \Q2[4] ,
    \Q2[3] ,
    \Q2[2] ,
    \Q2[1] ,
    \Q2[0] }),
    .Q3({\Q3[7] ,
    \Q3[6] ,
    \Q3[5] ,
    \Q3[4] ,
    \Q3[3] ,
    \Q3[2] ,
    \Q3[1] ,
    \Q3[0] }),
    .Q4({\Q4[7] ,
    \Q4[6] ,
    \Q4[5] ,
    \Q4[4] ,
    \Q4[3] ,
    \Q4[2] ,
    \Q4[1] ,
    \Q4[0] }),
    .Q5({\Q5[7] ,
    \Q5[6] ,
    \Q5[5] ,
    \Q5[4] ,
    \Q5[3] ,
    \Q5[2] ,
    \Q5[1] ,
    \Q5[0] }),
    .Q6({\Q6[7] ,
    \Q6[6] ,
    \Q6[5] ,
    \Q6[4] ,
    \Q6[3] ,
    \Q6[2] ,
    \Q6[1] ,
    \Q6[0] }),
    .Q7({\Q7[7] ,
    \Q7[6] ,
    \Q7[5] ,
    \Q7[4] ,
    \Q7[3] ,
    \Q7[2] ,
    \Q7[1] ,
    \Q7[0] }),
    .WEN_all({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }),
    .bus_in({\rom_bus_out[7] ,
    \rom_bus_out[6] ,
    \rom_bus_out[5] ,
    \rom_bus_out[4] ,
    \rom_bus_out[3] ,
    \rom_bus_out[2] ,
    \rom_bus_out[1] ,
    \rom_bus_out[0] }),
    .bus_out({\ram_bus_in[7] ,
    \ram_bus_in[6] ,
    \ram_bus_in[5] ,
    \ram_bus_in[4] ,
    \ram_bus_in[3] ,
    \ram_bus_in[2] ,
    \ram_bus_in[1] ,
    \ram_bus_in[0] }),
    .requested_addr({\requested_addr[15] ,
    \requested_addr[14] ,
    \requested_addr[13] ,
    \requested_addr[12] ,
    \requested_addr[11] ,
    \requested_addr[10] ,
    \requested_addr[9] ,
    \requested_addr[8] ,
    \requested_addr[7] ,
    \requested_addr[6] ,
    \requested_addr[5] ,
    \requested_addr[4] ,
    \requested_addr[3] ,
    \requested_addr[2] ,
    \requested_addr[1] ,
    \requested_addr[0] }));
 gf180mcu_fd_io__in_c rst_n_pad (.DVDD(VDD),
    .DVSS(VSS),
    .PAD(rst_n_PAD),
    .PD(\const_zero[1] ),
    .PU(\const_zero[0] ),
    .VDD(VDD),
    .VSS(VSS),
    .Y(rst_n_PAD2CORE));
 serial_ports serial_ports (.RXD(RXD),
    .TXD(TXD),
    .VDD(VDD),
    .VSS(VSS),
    .bus_cyc(bus_cyc),
    .bus_we(bus_we_serial_ports),
    .clk_i(clk_PAD2CORE),
    .io_in(\bidir_PAD2CORE[37] ),
    .irq3(irq3),
    .rst(reset),
    .addr({\bus_addr[2] ,
    \bus_addr[1] ,
    \bus_addr[0] }),
    .data_in({\bus_data_out[7] ,
    \bus_data_out[6] ,
    \bus_data_out[5] ,
    \bus_data_out[4] ,
    \bus_data_out[3] ,
    \bus_data_out[2] ,
    \bus_data_out[1] ,
    \bus_data_out[0] }),
    .data_out({\bus_data_serial_ports[7] ,
    \bus_data_serial_ports[6] ,
    \bus_data_serial_ports[5] ,
    \bus_data_serial_ports[4] ,
    \bus_data_serial_ports[3] ,
    \bus_data_serial_ports[2] ,
    \bus_data_serial_ports[1] ,
    \bus_data_serial_ports[0] }),
    .io_cs({\bidir_CORE2PAD_CS[37] ,
    \bidir_CORE2PAD_CS[36] ,
    \bidir_CORE2PAD_CS[35] }),
    .io_ie({\bidir_CORE2PAD_IE[37] ,
    \bidir_CORE2PAD_IE[36] ,
    \bidir_CORE2PAD_IE[35] }),
    .io_oe({\bidir_CORE2PAD_OE[37] ,
    \bidir_CORE2PAD_OE[36] ,
    \bidir_CORE2PAD_OE[35] }),
    .io_out({\bidir_CORE2PAD[37] ,
    \bidir_CORE2PAD[36] ,
    \bidir_CORE2PAD[35] }),
    .io_pd({\bidir_CORE2PAD_PD[37] ,
    \bidir_CORE2PAD_PD[36] ,
    \bidir_CORE2PAD_PD[35] }),
    .io_pu({\bidir_CORE2PAD_PU[37] ,
    \bidir_CORE2PAD_PU[36] ,
    \bidir_CORE2PAD_PU[35] }),
    .io_sl({\bidir_CORE2PAD_SL[37] ,
    \bidir_CORE2PAD_SL[36] ,
    \bidir_CORE2PAD_SL[35] }));
 sid sid (.DAC_clk(DAC_clk),
    .DAC_dat_1(DAC_d1),
    .DAC_dat_2(DAC_d2),
    .DAC_le(DAC_le),
    .VDD(VDD),
    .VSS(VSS),
    .bus_cyc(bus_cyc),
    .bus_we(bus_we_sid),
    .clk(clk_PAD2CORE),
    .rst(reset),
    .addr({\bus_addr[5] ,
    \bus_addr[4] ,
    \bus_addr[3] ,
    \bus_addr[2] ,
    \bus_addr[1] ,
    \bus_addr[0] }),
    .bus_in({\bus_data_out[7] ,
    \bus_data_out[6] ,
    \bus_data_out[5] ,
    \bus_data_out[4] ,
    \bus_data_out[3] ,
    \bus_data_out[2] ,
    \bus_data_out[1] ,
    \bus_data_out[0] }),
    .bus_out({\bus_data_sid[7] ,
    \bus_data_sid[6] ,
    \bus_data_sid[5] ,
    \bus_data_sid[4] ,
    \bus_data_sid[3] ,
    \bus_data_sid[2] ,
    \bus_data_sid[1] ,
    \bus_data_sid[0] }));
 gf180_ram_512x8_wrapper_as2650 sram0 (.CEN(CEN_all),
    .CLK(clk_PAD2CORE),
    .GWEN(GWEN_0),
    .VDD(VDD),
    .VSS(VSS),
    .A({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q({\Q0[7] ,
    \Q0[6] ,
    \Q0[5] ,
    \Q0[4] ,
    \Q0[3] ,
    \Q0[2] ,
    \Q0[1] ,
    \Q0[0] }),
    .WEN({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }));
 gf180_ram_512x8_wrapper_as2650 sram1 (.CEN(CEN_all),
    .CLK(clk_PAD2CORE),
    .GWEN(GWEN_1),
    .VDD(VDD),
    .VSS(VSS),
    .A({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q({\Q1[7] ,
    \Q1[6] ,
    \Q1[5] ,
    \Q1[4] ,
    \Q1[3] ,
    \Q1[2] ,
    \Q1[1] ,
    \Q1[0] }),
    .WEN({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }));
 gf180_ram_512x8_wrapper_as2650 sram2 (.CEN(CEN_all),
    .CLK(clk_PAD2CORE),
    .GWEN(GWEN_2),
    .VDD(VDD),
    .VSS(VSS),
    .A({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q({\Q2[7] ,
    \Q2[6] ,
    \Q2[5] ,
    \Q2[4] ,
    \Q2[3] ,
    \Q2[2] ,
    \Q2[1] ,
    \Q2[0] }),
    .WEN({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }));
 gf180_ram_512x8_wrapper_as2650 sram3 (.CEN(CEN_all),
    .CLK(clk_PAD2CORE),
    .GWEN(GWEN_3),
    .VDD(VDD),
    .VSS(VSS),
    .A({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q({\Q3[7] ,
    \Q3[6] ,
    \Q3[5] ,
    \Q3[4] ,
    \Q3[3] ,
    \Q3[2] ,
    \Q3[1] ,
    \Q3[0] }),
    .WEN({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }));
 gf180_ram_512x8_wrapper_as2650 sram4 (.CEN(CEN_all),
    .CLK(clk_PAD2CORE),
    .GWEN(GWEN_4),
    .VDD(VDD),
    .VSS(VSS),
    .A({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q({\Q4[7] ,
    \Q4[6] ,
    \Q4[5] ,
    \Q4[4] ,
    \Q4[3] ,
    \Q4[2] ,
    \Q4[1] ,
    \Q4[0] }),
    .WEN({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }));
 gf180_ram_512x8_wrapper_as2650 sram5 (.CEN(CEN_all),
    .CLK(clk_PAD2CORE),
    .GWEN(GWEN_5),
    .VDD(VDD),
    .VSS(VSS),
    .A({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q({\Q5[7] ,
    \Q5[6] ,
    \Q5[5] ,
    \Q5[4] ,
    \Q5[3] ,
    \Q5[2] ,
    \Q5[1] ,
    \Q5[0] }),
    .WEN({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }));
 gf180_ram_512x8_wrapper_as2650 sram6 (.CEN(CEN_all),
    .CLK(clk_PAD2CORE),
    .GWEN(GWEN_6),
    .VDD(VDD),
    .VSS(VSS),
    .A({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q({\Q6[7] ,
    \Q6[6] ,
    \Q6[5] ,
    \Q6[4] ,
    \Q6[3] ,
    \Q6[2] ,
    \Q6[1] ,
    \Q6[0] }),
    .WEN({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }));
 gf180_ram_512x8_wrapper_as2650 sram7 (.CEN(CEN_all),
    .CLK(clk_PAD2CORE),
    .GWEN(GWEN_7),
    .VDD(VDD),
    .VSS(VSS),
    .A({\A_all[8] ,
    \A_all[7] ,
    \A_all[6] ,
    \A_all[5] ,
    \A_all[4] ,
    \A_all[3] ,
    \A_all[2] ,
    \A_all[1] ,
    \A_all[0] }),
    .D({\D_all[7] ,
    \D_all[6] ,
    \D_all[5] ,
    \D_all[4] ,
    \D_all[3] ,
    \D_all[2] ,
    \D_all[1] ,
    \D_all[0] }),
    .Q({\Q7[7] ,
    \Q7[6] ,
    \Q7[5] ,
    \Q7[4] ,
    \Q7[3] ,
    \Q7[2] ,
    \Q7[1] ,
    \Q7[0] }),
    .WEN({\WEN_all[7] ,
    \WEN_all[6] ,
    \WEN_all[5] ,
    \WEN_all[4] ,
    \WEN_all[3] ,
    \WEN_all[2] ,
    \WEN_all[1] ,
    \WEN_all[0] }));
 timers timers (.VDD(VDD),
    .VSS(VSS),
    .bus_cyc(bus_cyc),
    .bus_we(bus_we_timers),
    .clk_i(clk_PAD2CORE),
    .irq1(irq1),
    .irq2(irq2),
    .irq5(irq5),
    .pwm0(pwm0),
    .pwm1(pwm1),
    .pwm2(pwm2),
    .rst(reset),
    .tmr0_clk(tmr0_clk),
    .tmr0_o(tmr0_o),
    .tmr1_clk(tmr1_clk),
    .tmr1_o(tmr1_o),
    .addr({\bus_addr[5] ,
    \bus_addr[4] ,
    \bus_addr[3] ,
    \bus_addr[2] ,
    \bus_addr[1] ,
    \bus_addr[0] }),
    .data_in({\bus_data_out[7] ,
    \bus_data_out[6] ,
    \bus_data_out[5] ,
    \bus_data_out[4] ,
    \bus_data_out[3] ,
    \bus_data_out[2] ,
    \bus_data_out[1] ,
    \bus_data_out[0] }),
    .data_out({\bus_data_timers[7] ,
    \bus_data_timers[6] ,
    \bus_data_timers[5] ,
    \bus_data_timers[4] ,
    \bus_data_timers[3] ,
    \bus_data_timers[2] ,
    \bus_data_timers[1] ,
    \bus_data_timers[0] }));
 unused unused (.VDD(VDD),
    .VSS(VSS),
    .clk_i(clk_PAD2CORE),
    .rst(reset),
    .io_cs({\bidir_CORE2PAD_CS[53] ,
    \bidir_CORE2PAD_CS[52] ,
    \bidir_CORE2PAD_CS[51] ,
    \bidir_CORE2PAD_CS[50] ,
    \bidir_CORE2PAD_CS[49] ,
    \bidir_CORE2PAD_CS[48] ,
    \bidir_CORE2PAD_CS[47] ,
    \bidir_CORE2PAD_CS[46] ,
    \bidir_CORE2PAD_CS[45] ,
    \bidir_CORE2PAD_CS[44] ,
    \bidir_CORE2PAD_CS[43] ,
    \bidir_CORE2PAD_CS[42] ,
    \bidir_CORE2PAD_CS[41] ,
    \bidir_CORE2PAD_CS[40] ,
    \bidir_CORE2PAD_CS[39] ,
    \bidir_CORE2PAD_CS[38] }),
    .io_ie({\bidir_CORE2PAD_IE[53] ,
    \bidir_CORE2PAD_IE[52] ,
    \bidir_CORE2PAD_IE[51] ,
    \bidir_CORE2PAD_IE[50] ,
    \bidir_CORE2PAD_IE[49] ,
    \bidir_CORE2PAD_IE[48] ,
    \bidir_CORE2PAD_IE[47] ,
    \bidir_CORE2PAD_IE[46] ,
    \bidir_CORE2PAD_IE[45] ,
    \bidir_CORE2PAD_IE[44] ,
    \bidir_CORE2PAD_IE[43] ,
    \bidir_CORE2PAD_IE[42] ,
    \bidir_CORE2PAD_IE[41] ,
    \bidir_CORE2PAD_IE[40] ,
    \bidir_CORE2PAD_IE[39] ,
    \bidir_CORE2PAD_IE[38] }),
    .io_in({\bidir_PAD2CORE[53] ,
    \bidir_PAD2CORE[52] ,
    \bidir_PAD2CORE[51] ,
    \bidir_PAD2CORE[50] ,
    \bidir_PAD2CORE[49] ,
    \bidir_PAD2CORE[48] ,
    \bidir_PAD2CORE[47] ,
    \bidir_PAD2CORE[46] ,
    \bidir_PAD2CORE[45] ,
    \bidir_PAD2CORE[44] ,
    \bidir_PAD2CORE[43] ,
    \bidir_PAD2CORE[42] ,
    \bidir_PAD2CORE[41] ,
    \bidir_PAD2CORE[40] ,
    \bidir_PAD2CORE[39] ,
    \bidir_PAD2CORE[38] }),
    .io_oe({\bidir_CORE2PAD_OE[53] ,
    \bidir_CORE2PAD_OE[52] ,
    \bidir_CORE2PAD_OE[51] ,
    \bidir_CORE2PAD_OE[50] ,
    \bidir_CORE2PAD_OE[49] ,
    \bidir_CORE2PAD_OE[48] ,
    \bidir_CORE2PAD_OE[47] ,
    \bidir_CORE2PAD_OE[46] ,
    \bidir_CORE2PAD_OE[45] ,
    \bidir_CORE2PAD_OE[44] ,
    \bidir_CORE2PAD_OE[43] ,
    \bidir_CORE2PAD_OE[42] ,
    \bidir_CORE2PAD_OE[41] ,
    \bidir_CORE2PAD_OE[40] ,
    \bidir_CORE2PAD_OE[39] ,
    \bidir_CORE2PAD_OE[38] }),
    .io_out({\bidir_CORE2PAD[53] ,
    \bidir_CORE2PAD[52] ,
    \bidir_CORE2PAD[51] ,
    \bidir_CORE2PAD[50] ,
    \bidir_CORE2PAD[49] ,
    \bidir_CORE2PAD[48] ,
    \bidir_CORE2PAD[47] ,
    \bidir_CORE2PAD[46] ,
    \bidir_CORE2PAD[45] ,
    \bidir_CORE2PAD[44] ,
    \bidir_CORE2PAD[43] ,
    \bidir_CORE2PAD[42] ,
    \bidir_CORE2PAD[41] ,
    \bidir_CORE2PAD[40] ,
    \bidir_CORE2PAD[39] ,
    \bidir_CORE2PAD[38] }),
    .io_pd({\bidir_CORE2PAD_PD[53] ,
    \bidir_CORE2PAD_PD[52] ,
    \bidir_CORE2PAD_PD[51] ,
    \bidir_CORE2PAD_PD[50] ,
    \bidir_CORE2PAD_PD[49] ,
    \bidir_CORE2PAD_PD[48] ,
    \bidir_CORE2PAD_PD[47] ,
    \bidir_CORE2PAD_PD[46] ,
    \bidir_CORE2PAD_PD[45] ,
    \bidir_CORE2PAD_PD[44] ,
    \bidir_CORE2PAD_PD[43] ,
    \bidir_CORE2PAD_PD[42] ,
    \bidir_CORE2PAD_PD[41] ,
    \bidir_CORE2PAD_PD[40] ,
    \bidir_CORE2PAD_PD[39] ,
    \bidir_CORE2PAD_PD[38] }),
    .io_pu({\bidir_CORE2PAD_PU[53] ,
    \bidir_CORE2PAD_PU[52] ,
    \bidir_CORE2PAD_PU[51] ,
    \bidir_CORE2PAD_PU[50] ,
    \bidir_CORE2PAD_PU[49] ,
    \bidir_CORE2PAD_PU[48] ,
    \bidir_CORE2PAD_PU[47] ,
    \bidir_CORE2PAD_PU[46] ,
    \bidir_CORE2PAD_PU[45] ,
    \bidir_CORE2PAD_PU[44] ,
    \bidir_CORE2PAD_PU[43] ,
    \bidir_CORE2PAD_PU[42] ,
    \bidir_CORE2PAD_PU[41] ,
    \bidir_CORE2PAD_PU[40] ,
    \bidir_CORE2PAD_PU[39] ,
    \bidir_CORE2PAD_PU[38] }),
    .io_sl({\bidir_CORE2PAD_SL[53] ,
    \bidir_CORE2PAD_SL[52] ,
    \bidir_CORE2PAD_SL[51] ,
    \bidir_CORE2PAD_SL[50] ,
    \bidir_CORE2PAD_SL[49] ,
    \bidir_CORE2PAD_SL[48] ,
    \bidir_CORE2PAD_SL[47] ,
    \bidir_CORE2PAD_SL[46] ,
    \bidir_CORE2PAD_SL[45] ,
    \bidir_CORE2PAD_SL[44] ,
    \bidir_CORE2PAD_SL[43] ,
    \bidir_CORE2PAD_SL[42] ,
    \bidir_CORE2PAD_SL[41] ,
    \bidir_CORE2PAD_SL[40] ,
    \bidir_CORE2PAD_SL[39] ,
    \bidir_CORE2PAD_SL[38] }));
 gf180mcu_ws_ip__logo wafer_space_logo ();
 wrapped_as2650 wrapped_as2650 (.VDD(VDD),
    .VSS(VSS),
    .WEb_ram(WEb_ram),
    .boot_rom_en(boot_rom_en),
    .bus_cyc(bus_cyc),
    .bus_we_gpios(bus_we_gpios),
    .bus_we_serial_ports(bus_we_serial_ports),
    .bus_we_sid(bus_we_sid),
    .bus_we_timers(bus_we_timers),
    .clk_i(clk_PAD2CORE),
    .le_hi_act(le_hi_act),
    .le_lo_act(le_lo_act),
    .ram_enabled(ram_enabled),
    .reset_out(reset),
    .rst_n(rst_n_PAD2CORE),
    .bus_addr({\bus_addr[5] ,
    \bus_addr[4] ,
    \bus_addr[3] ,
    \bus_addr[2] ,
    \bus_addr[1] ,
    \bus_addr[0] }),
    .bus_data_out({\bus_data_out[7] ,
    \bus_data_out[6] ,
    \bus_data_out[5] ,
    \bus_data_out[4] ,
    \bus_data_out[3] ,
    \bus_data_out[2] ,
    \bus_data_out[1] ,
    \bus_data_out[0] }),
    .bus_in_gpios({\bus_data_gpios[7] ,
    \bus_data_gpios[6] ,
    \bus_data_gpios[5] ,
    \bus_data_gpios[4] ,
    \bus_data_gpios[3] ,
    \bus_data_gpios[2] ,
    \bus_data_gpios[1] ,
    \bus_data_gpios[0] }),
    .bus_in_serial_ports({\bus_data_serial_ports[7] ,
    \bus_data_serial_ports[6] ,
    \bus_data_serial_ports[5] ,
    \bus_data_serial_ports[4] ,
    \bus_data_serial_ports[3] ,
    \bus_data_serial_ports[2] ,
    \bus_data_serial_ports[1] ,
    \bus_data_serial_ports[0] }),
    .bus_in_sid({\bus_data_sid[7] ,
    \bus_data_sid[6] ,
    \bus_data_sid[5] ,
    \bus_data_sid[4] ,
    \bus_data_sid[3] ,
    \bus_data_sid[2] ,
    \bus_data_sid[1] ,
    \bus_data_sid[0] }),
    .bus_in_timers({\bus_data_timers[7] ,
    \bus_data_timers[6] ,
    \bus_data_timers[5] ,
    \bus_data_timers[4] ,
    \bus_data_timers[3] ,
    \bus_data_timers[2] ,
    \bus_data_timers[1] ,
    \bus_data_timers[0] }),
    .const_zero({\const_zero[3] ,
    \const_zero[2] ,
    \const_zero[1] ,
    \const_zero[0] }),
    .io_cs({\bidir_CORE2PAD_CS[18] ,
    \bidir_CORE2PAD_CS[17] ,
    \bidir_CORE2PAD_CS[16] ,
    \bidir_CORE2PAD_CS[15] ,
    \bidir_CORE2PAD_CS[14] ,
    \bidir_CORE2PAD_CS[13] ,
    \bidir_CORE2PAD_CS[12] ,
    \bidir_CORE2PAD_CS[11] ,
    \bidir_CORE2PAD_CS[10] ,
    \bidir_CORE2PAD_CS[9] ,
    \bidir_CORE2PAD_CS[8] ,
    \bidir_CORE2PAD_CS[7] ,
    \bidir_CORE2PAD_CS[6] ,
    \bidir_CORE2PAD_CS[5] ,
    \bidir_CORE2PAD_CS[4] ,
    \bidir_CORE2PAD_CS[3] ,
    \bidir_CORE2PAD_CS[2] ,
    \bidir_CORE2PAD_CS[1] ,
    \bidir_CORE2PAD_CS[0] }),
    .io_ie({\bidir_CORE2PAD_IE[18] ,
    \bidir_CORE2PAD_IE[17] ,
    \bidir_CORE2PAD_IE[16] ,
    \bidir_CORE2PAD_IE[15] ,
    \bidir_CORE2PAD_IE[14] ,
    \bidir_CORE2PAD_IE[13] ,
    \bidir_CORE2PAD_IE[12] ,
    \bidir_CORE2PAD_IE[11] ,
    \bidir_CORE2PAD_IE[10] ,
    \bidir_CORE2PAD_IE[9] ,
    \bidir_CORE2PAD_IE[8] ,
    \bidir_CORE2PAD_IE[7] ,
    \bidir_CORE2PAD_IE[6] ,
    \bidir_CORE2PAD_IE[5] ,
    \bidir_CORE2PAD_IE[4] ,
    \bidir_CORE2PAD_IE[3] ,
    \bidir_CORE2PAD_IE[2] ,
    \bidir_CORE2PAD_IE[1] ,
    \bidir_CORE2PAD_IE[0] }),
    .io_in({\bidir_PAD2CORE[18] ,
    \bidir_PAD2CORE[17] ,
    \bidir_PAD2CORE[16] ,
    \bidir_PAD2CORE[15] ,
    \bidir_PAD2CORE[14] ,
    \bidir_PAD2CORE[13] ,
    \bidir_PAD2CORE[12] ,
    \bidir_PAD2CORE[11] ,
    \bidir_PAD2CORE[10] ,
    \bidir_PAD2CORE[9] ,
    \bidir_PAD2CORE[8] ,
    \bidir_PAD2CORE[7] ,
    \bidir_PAD2CORE[6] ,
    \bidir_PAD2CORE[5] ,
    \bidir_PAD2CORE[4] ,
    \bidir_PAD2CORE[3] ,
    \bidir_PAD2CORE[2] ,
    \bidir_PAD2CORE[1] ,
    \bidir_PAD2CORE[0] }),
    .io_oe({\bidir_CORE2PAD_OE[18] ,
    \bidir_CORE2PAD_OE[17] ,
    \bidir_CORE2PAD_OE[16] ,
    \bidir_CORE2PAD_OE[15] ,
    \bidir_CORE2PAD_OE[14] ,
    \bidir_CORE2PAD_OE[13] ,
    \bidir_CORE2PAD_OE[12] ,
    \bidir_CORE2PAD_OE[11] ,
    \bidir_CORE2PAD_OE[10] ,
    \bidir_CORE2PAD_OE[9] ,
    \bidir_CORE2PAD_OE[8] ,
    \bidir_CORE2PAD_OE[7] ,
    \bidir_CORE2PAD_OE[6] ,
    \bidir_CORE2PAD_OE[5] ,
    \bidir_CORE2PAD_OE[4] ,
    \bidir_CORE2PAD_OE[3] ,
    \bidir_CORE2PAD_OE[2] ,
    \bidir_CORE2PAD_OE[1] ,
    \bidir_CORE2PAD_OE[0] }),
    .io_out({\bidir_CORE2PAD[18] ,
    \bidir_CORE2PAD[17] ,
    \bidir_CORE2PAD[16] ,
    \bidir_CORE2PAD[15] ,
    \bidir_CORE2PAD[14] ,
    \bidir_CORE2PAD[13] ,
    \bidir_CORE2PAD[12] ,
    \bidir_CORE2PAD[11] ,
    \bidir_CORE2PAD[10] ,
    \bidir_CORE2PAD[9] ,
    \bidir_CORE2PAD[8] ,
    \bidir_CORE2PAD[7] ,
    \bidir_CORE2PAD[6] ,
    \bidir_CORE2PAD[5] ,
    \bidir_CORE2PAD[4] ,
    \bidir_CORE2PAD[3] ,
    \bidir_CORE2PAD[2] ,
    \bidir_CORE2PAD[1] ,
    \bidir_CORE2PAD[0] }),
    .io_pd({\bidir_CORE2PAD_PD[18] ,
    \bidir_CORE2PAD_PD[17] ,
    \bidir_CORE2PAD_PD[16] ,
    \bidir_CORE2PAD_PD[15] ,
    \bidir_CORE2PAD_PD[14] ,
    \bidir_CORE2PAD_PD[13] ,
    \bidir_CORE2PAD_PD[12] ,
    \bidir_CORE2PAD_PD[11] ,
    \bidir_CORE2PAD_PD[10] ,
    \bidir_CORE2PAD_PD[9] ,
    \bidir_CORE2PAD_PD[8] ,
    \bidir_CORE2PAD_PD[7] ,
    \bidir_CORE2PAD_PD[6] ,
    \bidir_CORE2PAD_PD[5] ,
    \bidir_CORE2PAD_PD[4] ,
    \bidir_CORE2PAD_PD[3] ,
    \bidir_CORE2PAD_PD[2] ,
    \bidir_CORE2PAD_PD[1] ,
    \bidir_CORE2PAD_PD[0] }),
    .io_pu({\bidir_CORE2PAD_PU[18] ,
    \bidir_CORE2PAD_PU[17] ,
    \bidir_CORE2PAD_PU[16] ,
    \bidir_CORE2PAD_PU[15] ,
    \bidir_CORE2PAD_PU[14] ,
    \bidir_CORE2PAD_PU[13] ,
    \bidir_CORE2PAD_PU[12] ,
    \bidir_CORE2PAD_PU[11] ,
    \bidir_CORE2PAD_PU[10] ,
    \bidir_CORE2PAD_PU[9] ,
    \bidir_CORE2PAD_PU[8] ,
    \bidir_CORE2PAD_PU[7] ,
    \bidir_CORE2PAD_PU[6] ,
    \bidir_CORE2PAD_PU[5] ,
    \bidir_CORE2PAD_PU[4] ,
    \bidir_CORE2PAD_PU[3] ,
    \bidir_CORE2PAD_PU[2] ,
    \bidir_CORE2PAD_PU[1] ,
    \bidir_CORE2PAD_PU[0] }),
    .io_sl({\bidir_CORE2PAD_SL[18] ,
    \bidir_CORE2PAD_SL[17] ,
    \bidir_CORE2PAD_SL[16] ,
    \bidir_CORE2PAD_SL[15] ,
    \bidir_CORE2PAD_SL[14] ,
    \bidir_CORE2PAD_SL[13] ,
    \bidir_CORE2PAD_SL[12] ,
    \bidir_CORE2PAD_SL[11] ,
    \bidir_CORE2PAD_SL[10] ,
    \bidir_CORE2PAD_SL[9] ,
    \bidir_CORE2PAD_SL[8] ,
    \bidir_CORE2PAD_SL[7] ,
    \bidir_CORE2PAD_SL[6] ,
    \bidir_CORE2PAD_SL[5] ,
    \bidir_CORE2PAD_SL[4] ,
    \bidir_CORE2PAD_SL[3] ,
    \bidir_CORE2PAD_SL[2] ,
    \bidir_CORE2PAD_SL[1] ,
    \bidir_CORE2PAD_SL[0] }),
    .irqs({irq7,
    irq6,
    irq5,
    irq3,
    irq2,
    irq1,
    irq0}),
    .last_addr({\last_addr[15] ,
    \last_addr[14] ,
    \last_addr[13] ,
    \last_addr[12] ,
    \last_addr[11] ,
    \last_addr[10] ,
    \last_addr[9] ,
    \last_addr[8] ,
    \last_addr[7] ,
    \last_addr[6] ,
    \last_addr[5] ,
    \last_addr[4] ,
    \last_addr[3] ,
    \last_addr[2] ,
    \last_addr[1] ,
    \last_addr[0] }),
    .ram_bus_in({\ram_bus_in[7] ,
    \ram_bus_in[6] ,
    \ram_bus_in[5] ,
    \ram_bus_in[4] ,
    \ram_bus_in[3] ,
    \ram_bus_in[2] ,
    \ram_bus_in[1] ,
    \ram_bus_in[0] }),
    .requested_addr({\requested_addr[15] ,
    \requested_addr[14] ,
    \requested_addr[13] ,
    \requested_addr[12] ,
    \requested_addr[11] ,
    \requested_addr[10] ,
    \requested_addr[9] ,
    \requested_addr[8] ,
    \requested_addr[7] ,
    \requested_addr[6] ,
    \requested_addr[5] ,
    \requested_addr[4] ,
    \requested_addr[3] ,
    \requested_addr[2] ,
    \requested_addr[1] ,
    \requested_addr[0] }),
    .rom_bus_in({\rom_bus_in[7] ,
    \rom_bus_in[6] ,
    \rom_bus_in[5] ,
    \rom_bus_in[4] ,
    \rom_bus_in[3] ,
    \rom_bus_in[2] ,
    \rom_bus_in[1] ,
    \rom_bus_in[0] }),
    .rom_bus_out({\rom_bus_out[7] ,
    \rom_bus_out[6] ,
    \rom_bus_out[5] ,
    \rom_bus_out[4] ,
    \rom_bus_out[3] ,
    \rom_bus_out[2] ,
    \rom_bus_out[1] ,
    \rom_bus_out[0] }));
 gf180mcu_fd_io__cor IO_CORNER_NORTH_WEST_INST (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__cor IO_CORNER_NORTH_EAST_INST (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__cor IO_CORNER_SOUTH_WEST_INST (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__cor IO_CORNER_SOUTH_EAST_INST (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_0_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_0_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_NORTH_0_1050 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_NORTH_0_1060 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_0_1070 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_0_1071 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_0_1072 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_0_1073 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_0_1074 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_1_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_1_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_2_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_2_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_3_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_3_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_4_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_4_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_5_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_5_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_6_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_6_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_7_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_7_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_8_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_8_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_9_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_9_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_10_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_10_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_11_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_11_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_12_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_12_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_13_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_13_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_14_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_14_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_15_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_15_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_16_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_16_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_NORTH_17_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_NORTH_17_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_NORTH_17_1050 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_NORTH_17_1060 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_17_1070 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_17_1071 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_17_1072 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_17_1073 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_NORTH_17_1074 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_0_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_0_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_SOUTH_0_1050 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_SOUTH_0_1060 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_0_1070 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_0_1071 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_0_1072 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_0_1073 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_0_1074 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_1_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_1_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_2_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_2_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_3_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_3_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_4_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_4_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_5_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_5_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_6_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_6_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_7_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_7_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_8_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_8_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_9_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_9_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_10_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_10_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_11_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_11_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_12_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_12_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_13_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_13_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_14_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_14_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_15_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_15_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_16_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_16_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_SOUTH_17_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_SOUTH_17_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_SOUTH_17_1050 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_SOUTH_17_1060 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_17_1070 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_17_1071 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_17_1072 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_17_1073 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fillnc IO_FILL_IO_SOUTH_17_1074 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_0_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_0_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_0_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_0_1360 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_0_1370 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_1_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_1_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_1_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_2_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_2_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_2_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_3_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_3_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_3_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_4_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_4_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_4_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_5_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_5_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_5_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_6_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_6_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_6_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_7_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_7_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_7_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_8_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_8_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_8_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_9_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_9_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_9_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_10_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_10_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_10_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_11_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_11_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_11_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_12_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_12_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_12_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_13_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_13_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_13_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_14_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_14_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_14_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_15_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_15_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_15_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_16_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_16_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_16_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_17_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_17_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_17_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_18_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_18_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_18_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_19_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_19_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_19_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_WEST_20_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_WEST_20_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_20_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_20_1360 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_WEST_20_1370 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_0_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_0_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_0_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_0_1360 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_0_1370 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_1_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_1_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_1_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_2_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_2_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_2_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_3_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_3_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_3_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_4_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_4_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_4_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_5_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_5_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_5_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_6_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_6_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_6_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_7_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_7_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_7_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_8_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_8_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_8_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_9_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_9_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_9_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_10_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_10_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_10_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_11_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_11_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_11_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_12_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_12_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_12_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_13_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_13_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_13_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_14_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_14_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_14_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_15_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_15_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_15_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_16_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_16_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_16_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_17_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_17_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_17_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_18_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_18_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_18_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_19_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_19_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_19_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_0 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_400 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_500 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_600 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_700 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_800 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_900 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_1000 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_1100 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill10 IO_FILL_IO_EAST_20_1200 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill5 IO_FILL_IO_EAST_20_1300 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_20_1350 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_20_1360 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_io__fill1 IO_FILL_IO_EAST_20_1370 (.DVDD(VDD),
    .DVSS(VSS),
    .VDD(VDD),
    .VSS(VSS));
endmodule
